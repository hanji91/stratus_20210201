/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:40:51 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755;
wire N5123,N5130,N5137,N5144,N5151,N5158,N5165 
	,N5172,N5179,N5186,N5193,N5200,N5207,N5214,N5221 
	,N5228,N5235,N5242,N5249,N5256,N5263,N5270,N5334 
	,N5336,N5572,N5585,N5587,N5611,N5613,N5676,N5683 
	,N5690,N5697,N5704,N5711,N5718,N5725,N5732,N5739 
	,N5746,N5753,N5760,N5767,N5774,N5781,N5788,N5795 
	,N5802,N5809,N5816,N5823,N5912,N5917,N5928,N5937 
	,N5946,N5955,N5964,N5973,N5982,N5991,N6000,N6153 
	,N6166,N6168,N6277,N6282,N6313,N6343,N6353,N6367 
	,N6369,N6400,N6419,N6425,N6427,N6451,N6456,N6458 
	,N6466,N6468,N6473,N6480,N6482,N6489,N6491,N6498 
	,N6507,N6509,N6516,N6525,N6527,N6534,N6543,N6545 
	,N6561,N6563,N6570,N6579,N6581,N6595,N6597,N6619 
	,N6649,N6688,N6737,N6794,N6851,N6909,N6967,N7025 
	,N7083,N7141,N7643,N7753,N7767,N7769,N7796,N7902 
	,N8095,N8097,N8099,N8182,N8198,N8261,N8556,N8564 
	,N8572,N8580,N8588,N8596,N8604,N8618,N8648,N8654 
	,N8663,N8670,N8677,N8684,N8691,N8699,N8707,N8715 
	,N8723,N8731,N8739,N8745,N8747,N8753,N8755,N8769 
	,N8779,N8781,N8787,N8797,N8799,N8805,N8815,N8817 
	,N8823,N8833,N8835,N8845,N8847,N8853,N8855,N8865 
	,N8867,N8873,N8875,N8885,N8887,N8893,N8895,N8905 
	,N8907,N8913,N8915,N8925,N8927,N8933,N8935,N8945 
	,N8947,N8953,N8955,N8965,N8967,N8977,N8981,N8983 
	,N9431,N9859;
EDFFHQX1 x_reg_L0_22__retimed_I4673 (.Q(N9431), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I4471 (.Q(N8983), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I4470 (.Q(N8981), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I4468 (.Q(N8977), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4463 (.Q(N8967), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4462 (.Q(N8965), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4458 (.Q(N8955), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4457 (.Q(N8953), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4455 (.Q(N8947), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4454 (.Q(N8945), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4450 (.Q(N8935), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4449 (.Q(N8933), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4447 (.Q(N8927), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4446 (.Q(N8925), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4442 (.Q(N8915), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4441 (.Q(N8913), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4439 (.Q(N8907), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4438 (.Q(N8905), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4434 (.Q(N8895), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4433 (.Q(N8893), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4431 (.Q(N8887), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4430 (.Q(N8885), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4426 (.Q(N8875), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4425 (.Q(N8873), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4423 (.Q(N8867), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4422 (.Q(N8865), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4418 (.Q(N8855), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4417 (.Q(N8853), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4415 (.Q(N8847), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4414 (.Q(N8845), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4410 (.Q(N8835), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4409 (.Q(N8833), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4405 (.Q(N8823), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4403 (.Q(N8817), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4402 (.Q(N8815), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4398 (.Q(N8805), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4396 (.Q(N8799), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4395 (.Q(N8797), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4391 (.Q(N8787), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4389 (.Q(N8781), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4388 (.Q(N8779), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4384 (.Q(N8769), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4379 (.Q(N8755), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4378 (.Q(N8753), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4377 (.Q(N8747), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4376 (.Q(N8745), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4375 (.Q(N8739), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4373 (.Q(N8731), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4371 (.Q(N8723), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4369 (.Q(N8715), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4367 (.Q(N8707), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4365 (.Q(N8699), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4363 (.Q(N8691), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4361 (.Q(N8684), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4359 (.Q(N8677), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4357 (.Q(N8670), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4355 (.Q(N8663), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4352 (.Q(N8654), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4351 (.Q(N8648), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4342 (.Q(N8618), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4338 (.Q(N8604), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4336 (.Q(N8596), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4334 (.Q(N8588), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4332 (.Q(N8580), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4330 (.Q(N8572), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4328 (.Q(N8564), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4326 (.Q(N8556), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4222 (.Q(N8261), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4197 (.Q(N8198), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4192 (.Q(N8182), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4173 (.Q(N8099), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4172 (.Q(N8097), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4171 (.Q(N8095), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4136 (.Q(N7902), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4112 (.Q(N7796), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4102 (.Q(N7769), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4101 (.Q(N7767), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I4095 (.Q(N7753), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I4061 (.Q(N7643), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3866 (.Q(N7141), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I3843 (.Q(N7083), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I3820 (.Q(N7025), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I3797 (.Q(N6967), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I3774 (.Q(N6909), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I3751 (.Q(N6851), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I3728 (.Q(N6794), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I3705 (.Q(N6737), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I3685 (.Q(N6688), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I3669 (.Q(N6649), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I3657 (.Q(N6619), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I3649 (.Q(N6597), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I3648 (.Q(N6595), .D(N6570), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_24__retimed_I3644 (.Q(N6581), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_24__retimed_I3643 (.Q(N6579), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3640 (.Q(N6570), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_25__retimed_I3638 (.Q(N6563), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_25__retimed_I3637 (.Q(N6561), .D(N6534), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_26__retimed_I3632 (.Q(N6545), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_26__retimed_I3631 (.Q(N6543), .D(N6516), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3628 (.Q(N6534), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_27__retimed_I3626 (.Q(N6527), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_27__retimed_I3625 (.Q(N6525), .D(N6498), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3622 (.Q(N6516), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_28__retimed_I3620 (.Q(N6509), .D(N6482), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_28__retimed_I3619 (.Q(N6507), .D(N6480), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3616 (.Q(N6498), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_29__retimed_I3614 (.Q(N6491), .D(N6458), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_29__retimed_I3613 (.Q(N6489), .D(N6456), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3611 (.Q(N6482), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3610 (.Q(N6480), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3608 (.Q(N6473), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_30__retimed_I3606 (.Q(N6468), .D(N6427), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_30__retimed_I3605 (.Q(N6466), .D(N6425), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3603 (.Q(N6458), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3602 (.Q(N6456), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3601 (.Q(N6451), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3591 (.Q(N6427), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3590 (.Q(N6425), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3589 (.Q(N6419), .D(N6353), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3582 (.Q(N6400), .D(N6343), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3569 (.Q(N6369), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3568 (.Q(N6367), .D(N6313), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3563 (.Q(N6353), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3560 (.Q(N6343), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3547 (.Q(N6313), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I3538 (.Q(N6282), .D(N5917), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I3536 (.Q(N6277), .D(N5912), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I3522 (.Q(N6168), .D(N5587), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I3521 (.Q(N6166), .D(N5585), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I3519 (.Q(N6153), .D(N5572), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I3461 (.Q(N6000), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I3457 (.Q(N5991), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I3453 (.Q(N5982), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I3449 (.Q(N5973), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I3445 (.Q(N5964), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I3441 (.Q(N5955), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I3437 (.Q(N5946), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I3433 (.Q(N5937), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I3429 (.Q(N5928), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_23__retimed_I3424 (.Q(N5917), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_7__retimed_I3422 (.Q(N5912), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I3413 (.Q(N5823), .D(N5270), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I3410 (.Q(N5816), .D(N5263), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I3407 (.Q(N5809), .D(N5256), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I3404 (.Q(N5802), .D(N5249), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I3401 (.Q(N5795), .D(N5242), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I3398 (.Q(N5788), .D(N5235), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I3395 (.Q(N5781), .D(N5228), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I3392 (.Q(N5774), .D(N5221), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I3389 (.Q(N5767), .D(N5214), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I3386 (.Q(N5760), .D(N5207), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I3383 (.Q(N5753), .D(N5200), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I3380 (.Q(N5746), .D(N5193), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I3377 (.Q(N5739), .D(N5186), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I3374 (.Q(N5732), .D(N5179), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I3371 (.Q(N5725), .D(N5172), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I3368 (.Q(N5718), .D(N5165), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I3365 (.Q(N5711), .D(N5158), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I3362 (.Q(N5704), .D(N5151), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I3359 (.Q(N5697), .D(N5144), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I3356 (.Q(N5690), .D(N5137), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I3353 (.Q(N5683), .D(N5130), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I3350 (.Q(N5676), .D(N5123), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_31__retimed_I3323 (.Q(N5613), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_31__retimed_I3322 (.Q(N5611), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_23__retimed_I3314 (.Q(N5587), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_23__retimed_I3313 (.Q(N5585), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I3311 (.Q(N5572), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_31__retimed_I3216 (.Q(N5336), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_31__retimed_I3215 (.Q(N5334), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I3188 (.Q(N5270), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_1__retimed_I3185 (.Q(N5263), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_2__retimed_I3182 (.Q(N5256), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_3__retimed_I3179 (.Q(N5249), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_4__retimed_I3176 (.Q(N5242), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_5__retimed_I3173 (.Q(N5235), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_6__retimed_I3170 (.Q(N5228), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_7__retimed_I3167 (.Q(N5221), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_8__retimed_I3164 (.Q(N5214), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_9__retimed_I3161 (.Q(N5207), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_10__retimed_I3158 (.Q(N5200), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_11__retimed_I3155 (.Q(N5193), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_12__retimed_I3152 (.Q(N5186), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_13__retimed_I3149 (.Q(N5179), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_14__retimed_I3146 (.Q(N5172), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_15__retimed_I3143 (.Q(N5165), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_16__retimed_I3140 (.Q(N5158), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_17__retimed_I3137 (.Q(N5151), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_18__retimed_I3134 (.Q(N5144), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_19__retimed_I3131 (.Q(N5137), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_20__retimed_I3128 (.Q(N5130), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I3125 (.Q(N5123), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21]), .E(bdw_enable), .CK(aclk));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149), .A(a_exp[7]), .B(a_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652), .A(a_man[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B(a_man[1]), .C(a_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134), .A(a_man[4]), .B(a_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157), .A(b_exp[7]), .B(b_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219), .A(b_man[4]), .B(b_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]));
OR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I46 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I47 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .A(b_exp[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I48 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .A(b_exp[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I49 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .A(b_exp[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I50 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .A(b_exp[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I51 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .A(b_exp[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I52 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558), .A(b_exp[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .A(b_exp[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .A(b_exp[0]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I56 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I57 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I58 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I59 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I60 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I61 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I62 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I66 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .B(a_exp[0]));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I67 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I68 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I69 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I70 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I71 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I72 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I73 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
OAI211X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950), .A(b_man[21]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633), .A(a_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642), .A(a_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459), .A(a_man[20]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241), .A(b_man[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386), .A(a_man[18]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387), .A(b_man[18]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369), .A(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371), .A(a_man[17]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378), .A(b_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384), .A(a_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378), .B(a_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264), .A(b_man[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427), .A(a_man[14]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428), .A(b_man[14]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410), .A(b_man[13]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412), .A(a_man[13]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419), .A(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425), .A(a_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419), .B(a_man[12]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287), .A(b_man[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468), .A(a_man[10]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469), .A(b_man[10]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451), .A(b_man[9]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453), .A(a_man[9]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461), .A(b_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466), .A(a_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461), .B(a_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310), .A(b_man[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319), .A(a_man[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323), .A(b_man[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346), .A(a_man[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333), .A(b_man[4]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351), .A(b_man[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344), .A(a_man[3]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975), .A(b_man[2]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975), .B(a_man[2]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980), .A(a_man[1]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I156 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I157 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986), .A(a_man[2]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I158 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I159 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981), .A(b_man[0]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I160 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977), .A(a_man[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I161 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972), .A0(b_man[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I162 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I163 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I166 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323), .B(a_man[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I167 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319), .B(b_man[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I168 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310), .B(a_man[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321));
AOI222X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I172 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430), .A(a_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298));
AOI222X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I176 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264), .B(a_man[15]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275));
AOI222X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I180 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241), .B(a_man[19]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252));
ACHCONX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I181 (.CON(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459), .B(b_man[20]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638), .B(b_man[22]));
AOI31X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575));
INVX12 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004), .A(b_man[20]), .B(a_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016), .A(b_man[19]), .B(a_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .B(a_exp[0]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .A(b_man[4]), .B(a_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .A(b_man[3]), .B(a_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .A(b_man[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .A(b_man[11]), .B(a_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .A(b_man[14]), .B(a_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .A(b_man[13]), .B(a_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835));
NOR4X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091));
NOR3X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .A(N8182), .B(N8198));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .A0N(N8965), .A1N(N8967), .B0(N8745), .B1(N8747));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .A0(N8739), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .B0(N8953), .B1(N8955));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .A0N(N8945), .A1N(N8947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .B1(N8731));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .A0(N8723), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .B0(N8933), .B1(N8935));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]));
AOI2BB2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .A0N(N8925), .A1N(N8927), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .B1(N8715));
OAI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .A0(N8707), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .B0(N8913), .B1(N8915));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .B(N8699));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .B(N8707));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .B(N8715));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .B(N8723));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .B(N8731));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .B(N8739));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .A(N8745), .B(N8747));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .A(N8753), .B(N8755));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I495 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664));
AOI2BB2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .A0N(N8905), .A1N(N8907), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .B1(N8699));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .A0(N8618), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .B0(N8893), .B1(N8895));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]));
AOI2BB2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .A0N(N8885), .A1N(N8887), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .B1(N8604));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .A0(N8596), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .B0(N8873), .B1(N8875));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]));
AOI2BB2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593), .A0N(N8865), .A1N(N8867), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .B1(N8588));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589), .A0(N8580), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593), .B0(N8853), .B1(N8855));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15]));
AOI2BB2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586), .A0N(N8845), .A1N(N8847), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589), .B1(N8572));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564), .A0(N8564), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586), .B0(N8833), .B1(N8835));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564), .B(N8556));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586), .B(N8564));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589), .B(N8572));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593), .B(N8580));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I527 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .B(N8588));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .B(N8596));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .B(N8604));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .B(N8618));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I535 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I549 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544), .A0(N8556), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564), .B0(N8823));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I550 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .A0(N8691), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544), .B0(N8815), .B1(N8817));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I552 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605), .A0(N8684), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .B0(N8805));
OAI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I553 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .A0(N8677), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605), .B0(N8797), .B1(N8799));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .B(N8670));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605), .B(N8677));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .B(N8684));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544), .B(N8691));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I564 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I566 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629), .A0(N8670), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .B0(N8787));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629), .B(N8663));
OAI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I572 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .A0(N8663), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629), .B0(N8779), .B1(N8781));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .B(N8648));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I579 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I582 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622), .A0(N8648), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .B0(N8769));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I583 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622), .B(N8654));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I584 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617), .A(N8654), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I585 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112), .A(N8095), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4617));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I586 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7112));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I589 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I590 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I591 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I601 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4750));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I607 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I608 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I610 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I612 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I614 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719), .A1(N8261), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I620 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I621 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I623 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I624 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4762), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4790));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I625 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I627 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I629 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I630 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I631 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4726), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4754));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I632 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4765), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4805));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I633 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4793));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I639 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780));
INVXL gen2_alt_A_I4887 (.Y(N9859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4716));
OAI2BB1X1 gen2_alt_A_I4888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .B0(N9859));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I641 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I644 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I645 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I647 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I648 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I649 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I650 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .A(N8198), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I661 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102), .A(N8182), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I673 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I680 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031), .A(N8198), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I690 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I691 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I692 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I693 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I694 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I695 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I696 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I697 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I698 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I699 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I700 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I701 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I706 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I713 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I714 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I715 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I716 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146), .A(N8182), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I735 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I750 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I751 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I752 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I758 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I761 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I762 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I768 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I770 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I771 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I773 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I774 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I779 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43), .A(N8097), .B(N8099), .S0(N8095));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I780 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I782 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I783 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548), .AN(a_sign), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565), .A(b_sign), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .A(rm[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .A(rm[1]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .C(rm[0]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I789 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .C(rm[0]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374), .A(N7902), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I794 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I795 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I796 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550), .A(N7902), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I797 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I798 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12550), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12592));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .B(rm[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5), .A(rm[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48), .A(a_sign), .B(b_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I804 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578), .A0(N7796), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12560), .B0(N7769));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I805 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636), .A(N7753), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12578));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I807 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54), .A(N7902), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I808 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639), .A0(N7767), .A1(N7769), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__54));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I809 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__53), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N636), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N639));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I810 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I811 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I812 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I813 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I814 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I815 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I816 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I817 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I818 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I819 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I820 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I821 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]), .A(N7643), .B(N8983));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I822 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]), .A(N7141), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I823 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]), .A(N7083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I824 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]), .A(N7025), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I825 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]), .A(N6967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I826 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]), .A(N6909), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I827 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]), .A(N6851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I828 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]), .A(N6794), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I829 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]), .A(N6737), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I830 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]), .A(N6688), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I831 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]), .A(N6649), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I832 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]), .A(N6619), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151), .A(N6473), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151), .B(N6451));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I840 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I848 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755), .B(N6419));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I851 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I852 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I853 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614), .A(N9431));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I856 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .A(N6597), .B(N6595), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I857 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .A(N6581), .B(N6579), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12123));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I858 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .A(N6563), .B(N6561), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12160));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I859 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]), .A(N6545), .B(N6543), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12194));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I860 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]), .A(N6527), .B(N6525), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12148));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I861 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .A(N6509), .B(N6507), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12184));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I862 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]), .A(N6491), .B(N6489), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12139));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I863 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]), .A(N6468), .B(N6466), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12174));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I864 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165), .A(N6400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I865 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125), .A(N6367), .B(N6369), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12165));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I866 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I867 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I868 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145), .A(N6400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12129));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I869 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12188), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12145));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I870 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12157), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12177));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I871 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12125), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12162));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I872 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__71));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
NOR2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .AN(N6153), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769), .A(rm[0]), .B(rm[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .B(N6277));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .A(N6153), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I885 (.Y(x[22]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[21]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[21]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I889 (.Y(x[21]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5676), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[20]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[20]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I892 (.Y(x[20]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5683), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I893 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[19]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I894 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I895 (.Y(x[19]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5690), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I896 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[18]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[18]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I897 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I898 (.Y(x[18]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5697), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I899 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[17]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I900 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I901 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I902 (.Y(x[17]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5704), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[16]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[16]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I905 (.Y(x[16]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5711), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I906 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[15]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[15]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I907 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I908 (.Y(x[15]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5718), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[14]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[14]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I911 (.Y(x[14]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5725), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[13]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I914 (.Y(x[13]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5732), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I915 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[12]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I916 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I918 (.Y(x[12]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5739), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[11]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[11]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I920 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I921 (.Y(x[11]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5746), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[10]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[10]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I923 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(N8981));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I924 (.Y(x[10]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5753), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I925 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[9]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(N8977));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I927 (.Y(x[9]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5760), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I928 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[8]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I929 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(N6000));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I930 (.Y(x[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5767), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5991));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I933 (.Y(x[7]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5774), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I935 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5982));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I936 (.Y(x[6]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5781), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I937 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I938 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5973));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I939 (.Y(x[5]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5788), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5964));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I942 (.Y(x[4]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5795), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5955));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I945 (.Y(x[3]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5802), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5946));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I948 (.Y(x[2]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5809), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5937));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I951 (.Y(x[1]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5816), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[0]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(N5928));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I954 (.Y(x[0]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N5823), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .A(N6168), .B(N6166), .C(N6153), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I957 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I958 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I959 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I960 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I961 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I962 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I963 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I964 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651), .A(N6282), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]), .A(N6166), .B(N6168), .C(N6153), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I967 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I968 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748), .A(a_sign), .B(b_sign));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952), .A0(a_sign), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_sign));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I974 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004), .A(N5611), .B(N5613), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I976 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[31]), .A(N5336), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004), .S0(N5334));
EDFFHQX1 x_reg_L1_31__I1040 (.Q(x[31]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[31]), .E(bdw_enable), .CK(aclk));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[29] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  v7DwSwDWqhw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



