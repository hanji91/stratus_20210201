/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:38:00 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
wire N5123,N5130,N5137,N5144,N5151,N5158,N5165 
	,N5172,N5179,N5186,N5193,N5200,N5207,N5214,N5221 
	,N5228,N5235,N5242,N5249,N5256,N5263,N5270,N5334 
	,N5336,N5572,N5588,N5590,N5614,N5616,N5700,N5705 
	,N5974,N6033,N6055,N6057,N6086,N6093,N6095,N6102 
	,N6138,N6147,N6523,N6777,N6784,N6860,N6930,N6937 
	,N6943,N6945,N6947,N6953,N7046,N7165,N7172,N7303 
	,N7323,N7343,N7350,N7357,N7364,N7371,N7379,N7421 
	,N7608,N7662,N7752,N7768,N7820,N7871,N7873,N7941 
	,N7946,N7955,N7962,N7969,N7976,N7983,N7990,N7997 
	,N8003,N8005,N8011,N8013,N8030,N8038,N8046,N8054 
	,N8062,N8070,N8078,N8086,N8148,N8522,N8527,N8533 
	,N8535,N8544,N9015,N9016,N9073,N9074,N9082,N9086 
	,N9088,N9100,N9101,N9115,N9117,N9121,N9123,N9125 
	,N9127,N9128,N9130,N9132,N9135,N9136,N9144,N9147 
	,N9149,N9151,N9156,N9158,N9161,N9163,N9168,N9172 
	,N9205,N9206,N9208,N9213,N9217,N9236,N9238,N9239 
	,N9261,N9265,N9267,N9269,N9273,N9294,N9298,N9303 
	,N9312,N9314,N9318,N9326,N9347,N9348,N9349,N9354 
	,N9355,N9361,N9373,N9377,N9381,N9385,N9387,N9391 
	,N9395,N9397,N9401,N9407,N9410,N9438,N9441,N9445 
	,N9448,N9459,N9464,N9469,N9474;
reg x_reg_22__retimed_I4614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4614_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3];
	end
assign N8544 = x_reg_22__retimed_I4614_QOUT;
reg x_reg_22__retimed_I4611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4611_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827;
	end
assign N8535 = x_reg_22__retimed_I4611_QOUT;
reg x_reg_22__retimed_I4610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4610_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831;
	end
assign N8533 = x_reg_22__retimed_I4610_QOUT;
reg x_reg_22__retimed_I4608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4608_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
	end
assign N8527 = x_reg_22__retimed_I4608_QOUT;
reg x_reg_22__retimed_I4606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4606_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4];
	end
assign N8522 = x_reg_22__retimed_I4606_QOUT;
reg x_reg_22__retimed_I4437_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4437_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N8148 = x_reg_22__retimed_I4437_QOUT;
reg x_reg_22__retimed_I4406_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4406_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679;
	end
assign N8086 = x_reg_22__retimed_I4406_QOUT;
reg x_reg_22__retimed_I4403_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4403_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609;
	end
assign N8078 = x_reg_22__retimed_I4403_QOUT;
reg x_reg_22__retimed_I4400_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4400_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687;
	end
assign N8070 = x_reg_22__retimed_I4400_QOUT;
reg x_reg_22__retimed_I4397_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4397_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618;
	end
assign N8062 = x_reg_22__retimed_I4397_QOUT;
reg x_reg_22__retimed_I4394_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4394_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695;
	end
assign N8054 = x_reg_22__retimed_I4394_QOUT;
reg x_reg_22__retimed_I4391_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4391_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626;
	end
assign N8046 = x_reg_22__retimed_I4391_QOUT;
reg x_reg_22__retimed_I4388_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4388_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704;
	end
assign N8038 = x_reg_22__retimed_I4388_QOUT;
reg x_reg_22__retimed_I4385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4385_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257;
	end
assign N8030 = x_reg_22__retimed_I4385_QOUT;
reg x_reg_22__retimed_I4380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4380_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722;
	end
assign N8013 = x_reg_22__retimed_I4380_QOUT;
reg x_reg_22__retimed_I4379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4379_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664;
	end
assign N8011 = x_reg_22__retimed_I4379_QOUT;
reg x_reg_22__retimed_I4378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4378_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636;
	end
assign N8005 = x_reg_22__retimed_I4378_QOUT;
reg x_reg_22__retimed_I4377_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4377_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659;
	end
assign N8003 = x_reg_22__retimed_I4377_QOUT;
reg x_reg_22__retimed_I4376_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4376_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700;
	end
assign N7997 = x_reg_22__retimed_I4376_QOUT;
reg x_reg_22__retimed_I4374_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4374_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620;
	end
assign N7990 = x_reg_22__retimed_I4374_QOUT;
reg x_reg_22__retimed_I4372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4372_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682;
	end
assign N7983 = x_reg_22__retimed_I4372_QOUT;
reg x_reg_22__retimed_I4370_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4370_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600;
	end
assign N7976 = x_reg_22__retimed_I4370_QOUT;
reg x_reg_22__retimed_I4368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4368_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665;
	end
assign N7969 = x_reg_22__retimed_I4368_QOUT;
reg x_reg_22__retimed_I4366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4366_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582;
	end
assign N7962 = x_reg_22__retimed_I4366_QOUT;
reg x_reg_22__retimed_I4364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4364_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644;
	end
assign N7955 = x_reg_22__retimed_I4364_QOUT;
reg x_reg_22__retimed_I4361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4361_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
	end
assign N7946 = x_reg_22__retimed_I4361_QOUT;
reg x_reg_22__retimed_I4360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4360_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677;
	end
assign N7941 = x_reg_22__retimed_I4360_QOUT;
reg x_reg_22__retimed_I4337_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4337_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894;
	end
assign N7873 = x_reg_22__retimed_I4337_QOUT;
reg x_reg_22__retimed_I4336_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4336_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914;
	end
assign N7871 = x_reg_22__retimed_I4336_QOUT;
reg x_reg_22__retimed_I4318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4318_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874;
	end
assign N7820 = x_reg_22__retimed_I4318_QOUT;
reg x_reg_22__retimed_I4300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4300_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840;
	end
assign N7768 = x_reg_22__retimed_I4300_QOUT;
reg x_reg_22__retimed_I4293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4293_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863;
	end
assign N7752 = x_reg_22__retimed_I4293_QOUT;
reg x_reg_22__retimed_I4272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4272_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896;
	end
assign N7662 = x_reg_22__retimed_I4272_QOUT;
reg x_reg_22__retimed_I4263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4263_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845;
	end
assign N7608 = x_reg_22__retimed_I4263_QOUT;
reg x_reg_22__retimed_I4235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4235_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486;
	end
assign N7421 = x_reg_22__retimed_I4235_QOUT;
reg x_reg_22__retimed_I4221_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4221_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N7379 = x_reg_22__retimed_I4221_QOUT;
reg x_reg_22__retimed_I4218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4218_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N7371 = x_reg_22__retimed_I4218_QOUT;
reg x_reg_22__retimed_I4215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N7364 = x_reg_22__retimed_I4215_QOUT;
reg x_reg_22__retimed_I4212_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4212_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N7357 = x_reg_22__retimed_I4212_QOUT;
reg x_reg_22__retimed_I4209_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4209_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N7350 = x_reg_22__retimed_I4209_QOUT;
reg x_reg_22__retimed_I4206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4206_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N7343 = x_reg_22__retimed_I4206_QOUT;
reg x_reg_22__retimed_I4198_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4198_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N7323 = x_reg_22__retimed_I4198_QOUT;
reg x_reg_22__retimed_I4191_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4191_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N7303 = x_reg_22__retimed_I4191_QOUT;
reg x_reg_22__retimed_I4157_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4157_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N7172 = x_reg_22__retimed_I4157_QOUT;
reg x_reg_22__retimed_I4154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4154_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N7165 = x_reg_22__retimed_I4154_QOUT;
reg x_reg_22__retimed_I4108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4108_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N7046 = x_reg_22__retimed_I4108_QOUT;
reg x_reg_22__retimed_I4071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N6953 = x_reg_22__retimed_I4071_QOUT;
reg x_reg_22__retimed_I4069_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4069_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N6947 = x_reg_22__retimed_I4069_QOUT;
reg x_reg_22__retimed_I4068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N6945 = x_reg_22__retimed_I4068_QOUT;
reg x_reg_22__retimed_I4067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4067_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N6943 = x_reg_22__retimed_I4067_QOUT;
reg x_reg_22__retimed_I4065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4065_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N6937 = x_reg_22__retimed_I4065_QOUT;
reg x_reg_22__retimed_I4062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4062_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N6930 = x_reg_22__retimed_I4062_QOUT;
reg x_reg_22__retimed_I4034_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4034_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N6860 = x_reg_22__retimed_I4034_QOUT;
reg x_reg_22__retimed_I4004_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4004_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N6784 = x_reg_22__retimed_I4004_QOUT;
reg x_reg_22__retimed_I4001_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4001_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N6777 = x_reg_22__retimed_I4001_QOUT;
reg x_reg_22__retimed_I3904_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3904_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N6523 = x_reg_22__retimed_I3904_QOUT;
reg x_reg_22__retimed_I3756_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3756_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N6147 = x_reg_22__retimed_I3756_QOUT;
reg x_reg_22__retimed_I3753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3753_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738;
	end
assign N6138 = x_reg_22__retimed_I3753_QOUT;
reg x_reg_22__retimed_I3741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3741_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
	end
assign N6102 = x_reg_22__retimed_I3741_QOUT;
reg x_reg_22__retimed_I3739_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3739_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439;
	end
assign N6095 = x_reg_22__retimed_I3739_QOUT;
reg x_reg_22__retimed_I3738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3738_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N6093 = x_reg_22__retimed_I3738_QOUT;
reg x_reg_22__retimed_I3736_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3736_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N6086 = x_reg_22__retimed_I3736_QOUT;
reg x_reg_22__retimed_I3727_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3727_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2];
	end
assign N6057 = x_reg_22__retimed_I3727_QOUT;
reg x_reg_22__retimed_I3726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3726_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N6055 = x_reg_22__retimed_I3726_QOUT;
reg x_reg_22__retimed_I3718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3718_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707;
	end
assign N6033 = x_reg_22__retimed_I3718_QOUT;
reg x_reg_22__retimed_I3695_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3695_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681;
	end
assign N5974 = x_reg_22__retimed_I3695_QOUT;
reg x_reg_23__retimed_I3594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3594_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N5705 = x_reg_23__retimed_I3594_QOUT;
reg x_reg_7__retimed_I3592_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3592_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912;
	end
assign N5700 = x_reg_7__retimed_I3592_QOUT;
reg x_reg_31__retimed_I3585_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3585_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N5616 = x_reg_31__retimed_I3585_QOUT;
reg x_reg_31__retimed_I3584_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3584_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5614 = x_reg_31__retimed_I3584_QOUT;
reg x_reg_23__retimed_I3576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3576_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5590 = x_reg_23__retimed_I3576_QOUT;
reg x_reg_23__retimed_I3575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3575_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5588 = x_reg_23__retimed_I3575_QOUT;
reg x_reg_22__retimed_I3572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3572_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5572 = x_reg_22__retimed_I3572_QOUT;
reg x_reg_31__retimed_I3477_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3477_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113;
	end
assign N5336 = x_reg_31__retimed_I3477_QOUT;
reg x_reg_31__retimed_I3476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3476_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122;
	end
assign N5334 = x_reg_31__retimed_I3476_QOUT;
reg x_reg_0__retimed_I3449_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3449_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5270 = x_reg_0__retimed_I3449_QOUT;
reg x_reg_1__retimed_I3446_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3446_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5263 = x_reg_1__retimed_I3446_QOUT;
reg x_reg_2__retimed_I3443_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3443_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5256 = x_reg_2__retimed_I3443_QOUT;
reg x_reg_3__retimed_I3440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3440_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5249 = x_reg_3__retimed_I3440_QOUT;
reg x_reg_4__retimed_I3437_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3437_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5242 = x_reg_4__retimed_I3437_QOUT;
reg x_reg_5__retimed_I3434_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3434_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5235 = x_reg_5__retimed_I3434_QOUT;
reg x_reg_6__retimed_I3431_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3431_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5228 = x_reg_6__retimed_I3431_QOUT;
reg x_reg_7__retimed_I3428_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3428_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5221 = x_reg_7__retimed_I3428_QOUT;
reg x_reg_8__retimed_I3425_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3425_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5214 = x_reg_8__retimed_I3425_QOUT;
reg x_reg_9__retimed_I3422_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3422_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5207 = x_reg_9__retimed_I3422_QOUT;
reg x_reg_10__retimed_I3419_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3419_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5200 = x_reg_10__retimed_I3419_QOUT;
reg x_reg_11__retimed_I3416_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3416_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5193 = x_reg_11__retimed_I3416_QOUT;
reg x_reg_12__retimed_I3413_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3413_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5186 = x_reg_12__retimed_I3413_QOUT;
reg x_reg_13__retimed_I3410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3410_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5179 = x_reg_13__retimed_I3410_QOUT;
reg x_reg_14__retimed_I3407_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3407_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5172 = x_reg_14__retimed_I3407_QOUT;
reg x_reg_15__retimed_I3404_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3404_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5165 = x_reg_15__retimed_I3404_QOUT;
reg x_reg_16__retimed_I3401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3401_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5158 = x_reg_16__retimed_I3401_QOUT;
reg x_reg_17__retimed_I3398_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3398_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5151 = x_reg_17__retimed_I3398_QOUT;
reg x_reg_18__retimed_I3395_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3395_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5144 = x_reg_18__retimed_I3395_QOUT;
reg x_reg_19__retimed_I3392_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3392_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5137 = x_reg_19__retimed_I3392_QOUT;
reg x_reg_20__retimed_I3389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3389_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5130 = x_reg_20__retimed_I3389_QOUT;
reg x_reg_21__retimed_I3386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3386_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5123 = x_reg_21__retimed_I3386_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123 = !(((a_man[0] | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168 = !(b_exp[0] & b_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202 = !((b_exp[7] & b_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056 = !(a_exp[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544 = !a_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426 = !(b_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479 = !(b_man[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410 = !a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530 = !(b_man[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433 = !(b_man[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485 = !(b_man[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537 = !(b_man[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489 = !a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496 = !(b_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550 = !(b_man[10] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451 = !(b_man[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453 = !a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439 = !(b_man[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492 = !(b_man[14] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542 = !(b_man[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446 = !(b_man[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503 = !(b_man[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525 = !a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404 = !(b_man[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455 = !(b_man[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547 = !a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506 = !(b_man[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408 = !(b_man[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460 = !(b_man[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527 = !(((a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475) | (b_man[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565} = {1'B0, a_exp[0]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 ^ a_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[11]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[13]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[4]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[4]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353)) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864);
assign N9459 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667 = !N9459;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[13]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[12]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[9]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign N9213 = N8003;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723 = (!N8086) | (N9213 & N8005);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] = (!N7997) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] = (!N8011) ^ N8013;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[17]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]);
assign N9205 = !(N8003 & N8005);
assign N9206 = !N7997;
assign N9217 = !((N9205 & N8086) | N9206);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699 = (!N8078) | (N7997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723);
assign N9208 = !N8078;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign N9361 = ((!N9217) & (!N9208)) | (!N7990);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597 = !(N8070 & N9361);
assign N9238 = (!N8062) | (N7983 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597);
assign N9464 = !N9238;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701 = !N9464;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578 = (!N8054) | (N7976 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578) ^ N7969;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597) ^ N7983;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699) ^ N7990;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign N9349 = !N8062;
assign N9347 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597 & N7983) | N9349);
assign N9355 = !N8054;
assign N9354 = !N7976;
assign N9348 = !(N9354 | N9347);
assign N9236 = !(N9355 | N9348);
assign N9239 = !N7969;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666 = (!N8046) | (N7969 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign N9448 = !N8046;
assign N9445 = !(N9239 | N9236);
assign N9438 = ((!N9445) & (!N9448)) | (!N7962);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672 = !(N8038 & N9438);
assign N9441 = !(N7955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594 = !(N8030 & N9441);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672) ^ N7955;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!N7962) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624 = !(N7941 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] = N7946 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900 = !(N7871 & N7873);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | N8148);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!N8003) ^ N8005;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701) ^ N7976;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24] = (!N7941) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907);
assign N9387 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | (!N8148));
assign N9397 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
assign N9407 = ((!N9387) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16])) | (!N9397);
assign N9373 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826) & (!N7820)) | (!N9407);
assign N9381 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
assign N9391 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
assign N9401 = ((!N9381) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20])) | (!N9391);
assign N9410 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
assign N9377 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
assign N9385 = ((!N9410) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24])) | (!N9377);
assign N9395 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855) & (!N9401)) | (!N9385);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 = !((N9373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892) | N9395);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841) & (!N7608)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[2]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729} = {1'B0, N6055} + {1'B0, N6057};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880 = !((N7768 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] = ((!N7662) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841) & (!N7752)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0];
assign N9073 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
assign N9074 = !N9073;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 = !(N8535 & N8533);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142;
assign N9261 = !N8533;
assign N9267 = !(N8535 | N9261);
assign N9269 = !(N8533 & (!N8535));
assign N9273 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892;
assign N9265 = !((N9267 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270 = (N9269 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842) | N9273;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174 = !(N9265 | N9273);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 & N7303;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign N9015 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177;
assign N9016 = !N9015;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]) | ((!N9016) & N6784);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285 = N7364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]) | ((!N9016) & N6930);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & N7165;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]) | ((!N9016) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & N7343;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]) | ((!N9016) & N8148);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214 = N7371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]) | ((!N9016) & N6937);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143 = N7379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & N7172);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & N7350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]) | ((!N9016) & N6523);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 & N7357;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]) | ((!N9016) & N6777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & N7172) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179) & N7379);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | ((!N9016) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146 = (N9016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]) | ((!N9016) & N7165);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & N8148) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & N7343);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & N6523) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & N7350);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & N6777) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N7357);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign N9298 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & N9298) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign N9314 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20] = !((N9314 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & N6784) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N7303);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] = !((N9314 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & N6930) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N7364);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & N9298) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & N6937) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N7371);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]);
assign N9318 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631 = N7421 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N7323) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280 = !(N6860 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N6953) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633 = N7046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269 = !(((N6943 | N6945) | N6947) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072;
assign N9469 = !N9318;
assign N9303 = !N9469;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596 = N9303 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign N9326 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]);
assign N9294 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]);
assign N9312 = !(N9318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543 = !((N9326 | N9294) | N9312);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 & a_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32) & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign N9086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & N9086) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213));
assign N9082 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & N9082) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248));
assign N9100 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543);
assign N9088 = N9100;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564 = !N9088;
assign N9101 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] = !(N9101 | N9100);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[3]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754} = {1'B0, N8544} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724} = {1'B0, N8522} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 & a_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433) & b_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 & a_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433) & b_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742 = !N8527;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446 = !N8527;
assign {N9158, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]} = {1'B0, N6147} + {1'B0, N9074} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]};
assign {N9125, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]} = {1'B0, N6138} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135} + {1'B0, N9158};
assign {N9151, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191} + {1'B0, N9125};
assign {N9117, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754} + {1'B0, N9151};
assign {N9144, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142} + {1'B0, N9117};
assign {N9168, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]} = {1'B0, N6102} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736} + {1'B0, N9144};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]} = {1'B0, N6093} + {1'B0, N6095} + {1'B0, N9168};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686} = {1'B0, N6086} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754 = !((N6055 & N6057) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642);
assign N9121 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]);
assign N9149 = !N9121;
assign N9115 = !((N9149 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]);
assign N9132 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]);
assign N9136 = !N9132;
assign N9163 = !(N9136 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign N9172 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683;
assign N9130 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62 = !(N6033 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754);
assign N9135 = !(N8527 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734);
assign N9128 = !(N5974 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]);
assign N9147 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62 | N9135);
assign N9156 = !(N9163 & N9115);
assign N9127 = !(N9172 & N9130);
assign N9161 = !((N9156 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686) | N9127);
assign N9123 = !(N9128 & N9147);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875 = !(N9123 | N9161);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 | (!N5572));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70 = N5700 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 = !(N5572 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5123);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5130);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5137);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5144);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5151);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5158);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5165);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5172);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5179);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5186);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5193);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5200);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5207);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5214);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5221);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5228);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5235);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5242);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5249);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5256);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5263);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[0]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N5270);
assign N9474 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] = !N9474;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869 = ((N5590 | N5588) | N5572) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651 = N5705 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0] = ((N5588 | N5590) | N5572) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] & N5616) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]) & N5614);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706);
assign x[31] = (N5334 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116) | ((!N5334) & N5336);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLXxTQrbrxA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



