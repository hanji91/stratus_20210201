`timescale 1ps / 1ps
module fix2float_Add_32Sx9S_32S_4_3(
          in2,
          in1,
          out1,
          clk
);
   input [31:0] in2;
   input [8:0] in1;
   output [31:0] out1;
   input clk;
wire add_23_2_n_0, add_23_2_n_1, add_23_2_n_2, add_23_2_n_3, add_23_2_n_4,
     add_23_2_n_5, add_23_2_n_6, add_23_2_n_7, add_23_2_n_8, add_23_2_n_9,
     add_23_2_n_10, add_23_2_n_11, add_23_2_n_12, add_23_2_n_13, add_23_2_n_14,
     add_23_2_n_15, add_23_2_n_16, add_23_2_n_17, add_23_2_n_18, add_23_2_n_19,
     add_23_2_n_20, add_23_2_n_21, add_23_2_n_22, add_23_2_n_23, add_23_2_n_24,
     add_23_2_n_25, add_23_2_n_26, add_23_2_n_27, add_23_2_n_28, add_23_2_n_29,
     add_23_2_n_30, add_23_2_n_31, add_23_2_n_32, add_23_2_n_33, add_23_2_n_34,
     add_23_2_n_35, add_23_2_n_36, add_23_2_n_37, add_23_2_n_38, add_23_2_n_39,
     add_23_2_n_40, add_23_2_n_41, add_23_2_n_42, add_23_2_n_43, add_23_2_n_44,
     add_23_2_n_45, add_23_2_n_46, add_23_2_n_47, add_23_2_n_48, add_23_2_n_49,
     add_23_2_n_50, add_23_2_n_51, add_23_2_n_52, add_23_2_n_53, add_23_2_n_54,
     add_23_2_n_55, add_23_2_n_56, add_23_2_n_57, add_23_2_n_58, add_23_2_n_59,
     add_23_2_n_60, add_23_2_n_61, add_23_2_n_62, add_23_2_n_63, add_23_2_n_64,
     add_23_2_n_65, add_23_2_n_66, add_23_2_n_67, add_23_2_n_68, add_23_2_n_69,
     add_23_2_n_70, add_23_2_n_71, add_23_2_n_72, add_23_2_n_74, add_23_2_n_75,
     add_23_2_n_76, add_23_2_n_77, add_23_2_n_78, add_23_2_n_79, add_23_2_n_80,
     add_23_2_n_81, add_23_2_n_82, add_23_2_n_83, add_23_2_n_84, add_23_2_n_85,
     add_23_2_n_86, add_23_2_n_87, add_23_2_n_88, add_23_2_n_89, add_23_2_n_90,
     add_23_2_n_91, add_23_2_n_92, add_23_2_n_93, add_23_2_n_95, add_23_2_n_96,
     add_23_2_n_97, add_23_2_n_98, add_23_2_n_99, add_23_2_n_100, add_23_2_n_103,
     add_23_2_n_107, add_23_2_n_111, add_23_2_n_112, add_23_2_n_113,
     add_23_2_n_114, add_23_2_n_115, add_23_2_n_116, add_23_2_n_117,
     add_23_2_n_118, add_23_2_n_122, add_23_2_n_128, add_23_2_n_129,
     add_23_2_n_131, add_23_2_n_132, add_23_2_n_134, add_23_2_n_135,
     add_23_2_n_136, add_23_2_n_139, add_23_2_n_140, add_23_2_n_141,
     add_23_2_n_144, add_23_2_n_145, add_23_2_n_146, add_23_2_n_147,
     add_23_2_n_148, add_23_2_n_152, add_23_2_n_153, add_23_2_n_154,
     add_23_2_n_156, add_23_2_n_157, add_23_2_n_158, add_23_2_n_162,
     add_23_2_n_163, add_23_2_n_164, add_23_2_n_168, add_23_2_n_169,
     add_23_2_n_170, add_23_2_n_173, add_23_2_n_174, add_23_2_n_175,
     add_23_2_n_179, add_23_2_n_180, add_23_2_n_183, add_23_2_n_186,
     add_23_2_n_187, add_23_2_n_190, add_23_2_n_191, n_18, n_20, n_22, n_23,
     n_25, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_39,
     n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_49, n_51, n_52, n_53, n_57,
     n_59, n_60, n_61, n_63, n_64, n_65, n_66, n_67, clk, n_110, n_111, n_114,
     n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, asc001_0_,
     asc001_1_, asc001_2_, asc001_3_, asc001_4_, asc001_5_, asc001_6_, asc001_7_,
     asc001_8_, asc001_9_, asc001_10_, asc001_11_, asc001_12_, asc001_13_,
     asc001_14_, asc001_15_, asc001_16_, asc001_17_, asc001_18_, asc001_19_,
     asc001_20_, asc001_21_, asc001_22_, asc001_23_, asc001_24_, asc001_25_,
     asc001_26_, asc001_27_, asc001_28_, asc001_29_, asc001_30_, asc001_31_;
assign {out1[31]} = asc001_31_;
assign {out1[30]} = asc001_30_;
assign {out1[29]} = asc001_29_;
assign {out1[28]} = asc001_28_;
assign {out1[27]} = asc001_27_;
assign {out1[26]} = asc001_26_;
assign {out1[25]} = asc001_25_;
assign {out1[24]} = asc001_24_;
assign {out1[23]} = asc001_23_;
assign {out1[22]} = asc001_22_;
assign {out1[21]} = asc001_21_;
assign {out1[20]} = asc001_20_;
assign {out1[19]} = asc001_19_;
assign {out1[18]} = asc001_18_;
assign {out1[17]} = asc001_17_;
assign {out1[15]} = asc001_15_;
assign {out1[14]} = asc001_14_;
assign {out1[13]} = asc001_13_;
 reg retime_s1_21_reg_reg_N30;
 always @(posedge clk)
         retime_s1_21_reg_reg_N30 <= add_23_2_n_93;
 assign n_39 = retime_s1_21_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         retime_s1_12_reg_reg_N30 <= add_23_2_n_2;
 assign n_51 = retime_s1_12_reg_reg_N30;
 reg retime_s1_35_reg_reg_N30;
 always @(posedge clk)
         retime_s1_35_reg_reg_N30 <= add_23_2_n_12;
 assign n_20 = retime_s1_35_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         retime_s1_13_reg_reg_N30 <= add_23_2_n_154;
 assign n_49 = retime_s1_13_reg_reg_N30;
 reg retime_s1_14_reg_reg_N30;
 always @(posedge clk)
         retime_s1_14_reg_reg_N30 <= add_23_2_n_89;
 assign n_46 = retime_s1_14_reg_reg_N30;
 reg retime_s1_15_reg_reg_N30;
 always @(posedge clk)
         retime_s1_15_reg_reg_N30 <= n_119;
 assign n_45 = retime_s1_15_reg_reg_N30;
 reg retime_s1_16_reg_reg_N30;
 always @(posedge clk)
         retime_s1_16_reg_reg_N30 <= add_23_2_n_61;
 assign n_44 = retime_s1_16_reg_reg_N30;
 reg retime_s1_17_reg_reg_N30;
 always @(posedge clk)
         retime_s1_17_reg_reg_N30 <= add_23_2_n_45;
 assign n_43 = retime_s1_17_reg_reg_N30;
 reg retime_s1_18_reg_reg_N30;
 always @(posedge clk)
         retime_s1_18_reg_reg_N30 <= {in2[26]};
 assign n_42 = retime_s1_18_reg_reg_N30;
 reg retime_s1_19_reg_reg_N30;
 always @(posedge clk)
         retime_s1_19_reg_reg_N30 <= add_23_2_n_42;
 assign n_41 = retime_s1_19_reg_reg_N30;
 reg retime_s1_27_reg_reg_N30;
 always @(posedge clk)
         retime_s1_27_reg_reg_N30 <= add_23_2_n_88;
 assign n_31 = retime_s1_27_reg_reg_N30;
 reg retime_s1_20_reg_reg_N30;
 always @(posedge clk)
         retime_s1_20_reg_reg_N30 <= add_23_2_n_75;
 assign n_40 = retime_s1_20_reg_reg_N30;
 reg out1_15_L0_reg_N30;
 always @(posedge clk)
         out1_15_L0_reg_N30 <= asc001_16_;
 assign {out1[16]} = out1_15_L0_reg_N30;
 reg retime_s1_22_reg_reg_N30;
 always @(posedge clk)
         retime_s1_22_reg_reg_N30 <= add_23_2_n_25;
 assign n_36 = retime_s1_22_reg_reg_N30;
 reg retime_s1_23_reg_reg_N30;
 always @(posedge clk)
         retime_s1_23_reg_reg_N30 <= add_23_2_n_91;
 assign n_35 = retime_s1_23_reg_reg_N30;
 reg retime_s1_24_reg_reg_N30;
 always @(posedge clk)
         retime_s1_24_reg_reg_N30 <= add_23_2_n_64;
 assign n_34 = retime_s1_24_reg_reg_N30;
 reg retime_s1_25_reg_reg_N30;
 always @(posedge clk)
         retime_s1_25_reg_reg_N30 <= add_23_2_n_20;
 assign n_33 = retime_s1_25_reg_reg_N30;
 reg retime_s1_26_reg_reg_N30;
 always @(posedge clk)
         retime_s1_26_reg_reg_N30 <= add_23_2_n_17;
 assign n_32 = retime_s1_26_reg_reg_N30;
 reg retime_s1_28_reg_reg_N30;
 always @(posedge clk)
         retime_s1_28_reg_reg_N30 <= add_23_2_n_13;
 assign n_30 = retime_s1_28_reg_reg_N30;
 reg retime_s1_29_reg_reg_N30;
 always @(posedge clk)
         retime_s1_29_reg_reg_N30 <= add_23_2_n_10;
 assign n_29 = retime_s1_29_reg_reg_N30;
 reg retime_s1_30_reg_reg_N30;
 always @(posedge clk)
         retime_s1_30_reg_reg_N30 <= add_23_2_n_96;
 assign n_28 = retime_s1_30_reg_reg_N30;
 reg retime_s1_31_reg_reg_N30;
 always @(posedge clk)
         retime_s1_31_reg_reg_N30 <= add_23_2_n_168;
 assign n_27 = retime_s1_31_reg_reg_N30;
 reg retime_s1_32_reg_reg_N30;
 always @(posedge clk)
         retime_s1_32_reg_reg_N30 <= add_23_2_n_0;
 assign n_25 = retime_s1_32_reg_reg_N30;
 reg retime_s1_33_reg_reg_N30;
 always @(posedge clk)
         retime_s1_33_reg_reg_N30 <= add_23_2_n_164;
 assign n_23 = retime_s1_33_reg_reg_N30;
 reg retime_s1_34_reg_reg_N30;
 always @(posedge clk)
         retime_s1_34_reg_reg_N30 <= add_23_2_n_153;
 assign n_22 = retime_s1_34_reg_reg_N30;
 reg out1_28_L0_reg_N30;
 always @(posedge clk)
         out1_28_L0_reg_N30 <= asc001_3_;
 assign {out1[3]} = out1_28_L0_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         retime_s1_11_reg_reg_N30 <= add_23_2_n_157;
 assign n_52 = retime_s1_11_reg_reg_N30;
 reg out1_19_L0_reg_N30;
 always @(posedge clk)
         out1_19_L0_reg_N30 <= asc001_12_;
 assign {out1[12]} = out1_19_L0_reg_N30;
 reg out1_20_L0_reg_N30;
 always @(posedge clk)
         out1_20_L0_reg_N30 <= asc001_11_;
 assign {out1[11]} = out1_20_L0_reg_N30;
 reg out1_21_L0_reg_N30;
 always @(posedge clk)
         out1_21_L0_reg_N30 <= asc001_10_;
 assign {out1[10]} = out1_21_L0_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         retime_s1_7_reg_reg_N30 <= add_23_2_n_163;
 assign n_60 = retime_s1_7_reg_reg_N30;
 reg out1_22_L0_reg_N30;
 always @(posedge clk)
         out1_22_L0_reg_N30 <= asc001_9_;
 assign {out1[9]} = out1_22_L0_reg_N30;
 reg out1_23_L0_reg_N30;
 always @(posedge clk)
         out1_23_L0_reg_N30 <= asc001_8_;
 assign {out1[8]} = out1_23_L0_reg_N30;
 reg out1_24_L0_reg_N30;
 always @(posedge clk)
         out1_24_L0_reg_N30 <= asc001_7_;
 assign {out1[7]} = out1_24_L0_reg_N30;
 reg out1_25_L0_reg_N30;
 always @(posedge clk)
         out1_25_L0_reg_N30 <= asc001_6_;
 assign {out1[6]} = out1_25_L0_reg_N30;
 reg out1_26_L0_reg_N30;
 always @(posedge clk)
         out1_26_L0_reg_N30 <= asc001_5_;
 assign {out1[5]} = out1_26_L0_reg_N30;
 reg out1_27_L0_reg_N30;
 always @(posedge clk)
         out1_27_L0_reg_N30 <= asc001_4_;
 assign {out1[4]} = out1_27_L0_reg_N30;
 reg retime_s1_36_reg_reg_N30;
 always @(posedge clk)
         retime_s1_36_reg_reg_N30 <= {in2[29]};
 assign n_18 = retime_s1_36_reg_reg_N30;
 reg out1_29_L0_reg_N30;
 always @(posedge clk)
         out1_29_L0_reg_N30 <= asc001_2_;
 assign {out1[2]} = out1_29_L0_reg_N30;
 reg out1_30_L0_reg_N30;
 always @(posedge clk)
         out1_30_L0_reg_N30 <= asc001_1_;
 assign {out1[1]} = out1_30_L0_reg_N30;
 reg out1_31_L0_reg_N30;
 always @(posedge clk)
         out1_31_L0_reg_N30 <= asc001_0_;
 assign {out1[0]} = out1_31_L0_reg_N30;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= {in2[30]};
 assign n_67 = retime_s1_1_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= n_114;
 assign n_65 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= add_23_2_n_59;
 assign n_64 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= add_23_2_n_69;
 assign n_63 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= add_23_2_n_58;
 assign n_61 = retime_s1_6_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         retime_s1_8_reg_reg_N30 <= add_23_2_n_156;
 assign n_59 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         retime_s1_9_reg_reg_N30 <= add_23_2_n_158;
 assign n_57 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         retime_s1_10_reg_reg_N30 <= add_23_2_n_66;
 assign n_53 = retime_s1_10_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= {in1[8]};
 assign n_66 = retime_s1_2_reg_reg_N30;
 assign asc001_31_ = ~(add_23_2_n_191 ^ n_61);
 assign add_23_2_n_191 = ((add_23_2_n_190 & n_67) | ((n_67 & n_66) | (n_66 & add_23_2_n_190)));
 assign asc001_30_ = (n_67 ^ (n_66 ^ add_23_2_n_190));
 assign add_23_2_n_190 = ~(add_23_2_n_56 & (add_23_2_n_187 | add_23_2_n_27));
 assign asc001_29_ = ~(add_23_2_n_186 ^ add_23_2_n_80);
 assign asc001_27_ = ~(add_23_2_n_183 ^ add_23_2_n_71);
 assign add_23_2_n_187 = ~(add_23_2_n_44 | (add_23_2_n_179 & n_33));
 assign add_23_2_n_186 = ~(n_43 & ~(add_23_2_n_179 & n_33));
 assign asc001_28_ = ~(add_23_2_n_179 ^ add_23_2_n_72);
 assign asc001_23_ = ~(add_23_2_n_180 ^ n_34);
 assign add_23_2_n_183 = ~(add_23_2_n_8 & (add_23_2_n_174 | add_23_2_n_40));
 assign asc001_26_ = ~(add_23_2_n_174 ^ add_23_2_n_83);
 assign asc001_25_ = ~(add_23_2_n_173 ^ n_63);
 assign add_23_2_n_180 = ~(n_30 & (add_23_2_n_170 | n_25));
 assign add_23_2_n_179 = ~(add_23_2_n_116 & (add_23_2_n_175 & (n_51 | add_23_2_n_8)));
 assign asc001_22_ = ~(add_23_2_n_170 ^ add_23_2_n_62);
 assign asc001_21_ = ~(add_23_2_n_169 ^ n_44);
 assign asc001_19_ = ~(n_27 ^ n_53);
 assign add_23_2_n_175 = ~(n_36 | (n_28 & (add_23_2_n_74 & n_60)));
 assign add_23_2_n_174 = ~(n_65 | (n_60 & n_28));
 assign add_23_2_n_173 = ~(n_20 & (add_23_2_n_162 | n_29));
 assign asc001_15_ = ~(n_23 ^ n_46);
 assign asc001_24_ = ~(n_60 ^ add_23_2_n_65);
 assign add_23_2_n_170 = ~(n_45 | (n_52 & n_40));
 assign add_23_2_n_169 = ~(n_32 & ~(n_52 & n_41));
 assign add_23_2_n_168 = ~(add_23_2_n_39 & (add_23_2_n_156 | add_23_2_n_7));
 assign asc001_18_ = ~(n_59 ^ n_39);
 assign asc001_17_ = ~(n_57 ^ n_35);
 assign asc001_20_ = ~(n_52 ^ add_23_2_n_60);
 assign add_23_2_n_164 = ~(add_23_2_n_16 & (add_23_2_n_154 | add_23_2_n_11));
 assign add_23_2_n_162 = ~n_60;
 assign add_23_2_n_163 = ~(n_111 & (add_23_2_n_147 | (add_23_2_n_112 | add_23_2_n_114)));
 assign asc001_14_ = ~(n_49 ^ n_31);
 assign asc001_13_ = ~(n_22 ^ n_64);
 assign asc001_11_ = ~(add_23_2_n_152 ^ add_23_2_n_63);
 assign add_23_2_n_158 = ~(add_23_2_n_15 & (add_23_2_n_147 | add_23_2_n_21));
 assign add_23_2_n_157 = ~(add_23_2_n_117 & (n_116 & (add_23_2_n_147 | add_23_2_n_112)));
 assign add_23_2_n_156 = ~(n_118 | (add_23_2_n_148 & add_23_2_n_95));
 assign asc001_16_ = ~(add_23_2_n_148 ^ add_23_2_n_90);
 assign add_23_2_n_154 = ~(n_120 | (add_23_2_n_146 & add_23_2_n_97));
 assign add_23_2_n_153 = ~(add_23_2_n_47 & ~(add_23_2_n_146 & add_23_2_n_43));
 assign add_23_2_n_152 = ~(add_23_2_n_30 & (add_23_2_n_144 | add_23_2_n_32));
 assign asc001_12_ = ~(add_23_2_n_146 ^ add_23_2_n_87);
 assign asc001_10_ = ~(add_23_2_n_144 ^ add_23_2_n_86);
 assign asc001_9_ = ~(add_23_2_n_145 ^ add_23_2_n_85);
 assign add_23_2_n_147 = ~add_23_2_n_148;
 assign add_23_2_n_148 = ~(n_110 & (add_23_2_n_139 | (add_23_2_n_111 | add_23_2_n_113)));
 assign add_23_2_n_146 = ~(add_23_2_n_115 & (n_117 & (add_23_2_n_139 | add_23_2_n_113)));
 assign add_23_2_n_145 = ~(add_23_2_n_5 & (add_23_2_n_139 | add_23_2_n_31));
 assign add_23_2_n_144 = ~(n_115 | (add_23_2_n_140 & add_23_2_n_100));
 assign asc001_8_ = ~(add_23_2_n_140 ^ add_23_2_n_67);
 assign asc001_7_ = ~(add_23_2_n_141 ^ add_23_2_n_84);
 assign add_23_2_n_141 = ~(add_23_2_n_46 & (add_23_2_n_135 | add_23_2_n_34));
 assign add_23_2_n_139 = ~add_23_2_n_140;
 assign add_23_2_n_140 = ~(add_23_2_n_118 & (add_23_2_n_136 & (add_23_2_n_3 | add_23_2_n_46)));
 assign asc001_6_ = ~(add_23_2_n_135 ^ add_23_2_n_68);
 assign asc001_5_ = ~(add_23_2_n_134 ^ add_23_2_n_70);
 assign add_23_2_n_136 = ~(add_23_2_n_51 | (add_23_2_n_132 & (add_23_2_n_78 & add_23_2_n_76)));
 assign add_23_2_n_135 = ~(add_23_2_n_103 | (add_23_2_n_132 & add_23_2_n_76));
 assign add_23_2_n_134 = ~(add_23_2_n_1 & (add_23_2_n_131 | add_23_2_n_41));
 assign asc001_4_ = ~(add_23_2_n_132 ^ add_23_2_n_82);
 assign add_23_2_n_131 = ~add_23_2_n_132;
 assign add_23_2_n_132 = ~(add_23_2_n_23 & (add_23_2_n_128 | add_23_2_n_24));
 assign asc001_3_ = ~(add_23_2_n_129 ^ add_23_2_n_81);
 assign add_23_2_n_129 = ~(add_23_2_n_19 & ~(add_23_2_n_122 & add_23_2_n_33));
 assign add_23_2_n_128 = ~(add_23_2_n_18 | (add_23_2_n_122 & add_23_2_n_33));
 assign asc001_2_ = ~(add_23_2_n_122 ^ add_23_2_n_92);
 assign add_23_2_n_122 = ((add_23_2_n_107 & {in2[1]}) | (({in2[1]} & {in1[1]}) | ({in1[1]} & add_23_2_n_107)));
 assign asc001_1_ = ({in2[1]} ^ ({in1[1]} ^ add_23_2_n_107));
 assign add_23_2_n_118 = ~(add_23_2_n_103 & add_23_2_n_78);
 assign add_23_2_n_116 = ~(n_65 & add_23_2_n_74);
 assign add_23_2_n_107 = ({in1[0]} & {in2[0]});
 assign asc001_0_ = ({in1[0]} ^ {in2[0]});
 assign add_23_2_n_114 = ~(add_23_2_n_75 & add_23_2_n_77);
 assign add_23_2_n_113 = ~(add_23_2_n_100 & add_23_2_n_98);
 assign add_23_2_n_112 = ~(add_23_2_n_95 & add_23_2_n_99);
 assign add_23_2_n_111 = ~(add_23_2_n_97 & add_23_2_n_79);
 assign add_23_2_n_103 = ~(add_23_2_n_48 & (add_23_2_n_36 | add_23_2_n_1));
 assign add_23_2_n_93 = ~(add_23_2_n_7 | ~add_23_2_n_39);
 assign add_23_2_n_92 = ~(add_23_2_n_33 & add_23_2_n_19);
 assign add_23_2_n_91 = ~(add_23_2_n_26 & ~add_23_2_n_14);
 assign add_23_2_n_90 = ~(add_23_2_n_15 & ~add_23_2_n_21);
 assign add_23_2_n_89 = ~(add_23_2_n_57 & ~add_23_2_n_37);
 assign add_23_2_n_100 = ~(add_23_2_n_31 | add_23_2_n_29);
 assign add_23_2_n_88 = ~(add_23_2_n_11 | ~add_23_2_n_16);
 assign add_23_2_n_87 = ~(add_23_2_n_43 & add_23_2_n_47);
 assign add_23_2_n_86 = ~(add_23_2_n_32 | ~add_23_2_n_30);
 assign add_23_2_n_85 = ~(add_23_2_n_52 & ~add_23_2_n_29);
 assign add_23_2_n_99 = ~(add_23_2_n_7 | add_23_2_n_6);
 assign add_23_2_n_98 = ~(add_23_2_n_32 | add_23_2_n_38);
 assign add_23_2_n_97 = ~(add_23_2_n_9 | ~add_23_2_n_43);
 assign add_23_2_n_84 = (add_23_2_n_3 | add_23_2_n_51);
 assign add_23_2_n_83 = ~(add_23_2_n_40 | ~add_23_2_n_8);
 assign add_23_2_n_82 = ~(add_23_2_n_1 & ~add_23_2_n_41);
 assign add_23_2_n_96 = ~(add_23_2_n_10 | add_23_2_n_4);
 assign add_23_2_n_95 = ~(add_23_2_n_21 | add_23_2_n_14);
 assign add_23_2_n_81 = ~(add_23_2_n_23 & ~add_23_2_n_24);
 assign add_23_2_n_80 = ~(add_23_2_n_56 & ~add_23_2_n_27);
 assign add_23_2_n_72 = ~(n_33 & n_43);
 assign add_23_2_n_79 = ~(add_23_2_n_11 | add_23_2_n_37);
 assign add_23_2_n_71 = (n_51 | n_36);
 assign add_23_2_n_70 = ~(add_23_2_n_48 & ~add_23_2_n_36);
 assign add_23_2_n_69 = ~(add_23_2_n_55 & ~add_23_2_n_4);
 assign add_23_2_n_68 = ~(add_23_2_n_34 | ~add_23_2_n_46);
 assign add_23_2_n_78 = ~(add_23_2_n_34 | add_23_2_n_3);
 assign add_23_2_n_67 = ~(add_23_2_n_5 & ~add_23_2_n_31);
 assign add_23_2_n_66 = ~(add_23_2_n_49 & ~add_23_2_n_6);
 assign add_23_2_n_77 = ~(add_23_2_n_0 | add_23_2_n_22);
 assign add_23_2_n_65 = ~(n_20 & ~n_29);
 assign add_23_2_n_64 = ~(add_23_2_n_53 & ~add_23_2_n_22);
 assign add_23_2_n_76 = ~(add_23_2_n_41 | add_23_2_n_36);
 assign add_23_2_n_63 = ~(add_23_2_n_28 & ~add_23_2_n_38);
 assign add_23_2_n_62 = ~(n_25 | ~n_30);
 assign add_23_2_n_61 = ~(add_23_2_n_50 & ~add_23_2_n_35);
 assign add_23_2_n_60 = ~(n_41 & n_32);
 assign add_23_2_n_75 = ~(add_23_2_n_35 | ~add_23_2_n_42);
 assign add_23_2_n_74 = ~(add_23_2_n_40 | n_51);
 assign add_23_2_n_59 = ~(add_23_2_n_54 & ~add_23_2_n_9);
 assign add_23_2_n_58 = ~({in1[8]} ^ {in2[31]});
 assign add_23_2_n_44 = ~n_43;
 assign add_23_2_n_57 = ~({in1[8]} & {in2[15]});
 assign add_23_2_n_56 = ~(n_66 & n_18);
 assign add_23_2_n_55 = ~({in1[8]} & {in2[25]});
 assign add_23_2_n_54 = ~({in1[8]} & {in2[13]});
 assign add_23_2_n_53 = ~({in1[8]} & {in2[23]});
 assign add_23_2_n_52 = ~({in1[8]} & {in2[9]});
 assign add_23_2_n_51 = ({in1[7]} & {in2[7]});
 assign add_23_2_n_50 = ~({in1[8]} & {in2[21]});
 assign add_23_2_n_49 = ~({in1[8]} & {in2[19]});
 assign add_23_2_n_48 = ~({in1[5]} & {in2[5]});
 assign add_23_2_n_47 = ~({in1[8]} & {in2[12]});
 assign add_23_2_n_46 = ~({in1[6]} & {in2[6]});
 assign add_23_2_n_45 = ~({in1[8]} & {in2[28]});
 assign add_23_2_n_43 = ({in1[8]} | {in2[12]});
 assign add_23_2_n_42 = ({in1[8]} | {in2[20]});
 assign add_23_2_n_41 = ~({in1[4]} | {in2[4]});
 assign add_23_2_n_40 = ~(n_66 | n_42);
 assign add_23_2_n_39 = ~({in1[8]} & {in2[18]});
 assign add_23_2_n_38 = ~({in1[8]} | {in2[11]});
 assign add_23_2_n_37 = ~({in1[8]} | {in2[15]});
 assign add_23_2_n_36 = ~({in1[5]} | {in2[5]});
 assign add_23_2_n_35 = ~({in1[8]} | {in2[21]});
 assign add_23_2_n_34 = ~({in1[6]} | {in2[6]});
 assign add_23_2_n_33 = ({in1[2]} | {in2[2]});
 assign add_23_2_n_32 = ~({in1[8]} | {in2[10]});
 assign add_23_2_n_31 = ~({in1[8]} | {in2[8]});
 assign add_23_2_n_30 = ~({in1[8]} & {in2[10]});
 assign add_23_2_n_29 = ~({in1[8]} | {in2[9]});
 assign add_23_2_n_18 = ~add_23_2_n_19;
 assign add_23_2_n_28 = ~({in1[8]} & {in2[11]});
 assign add_23_2_n_27 = ~(n_66 | n_18);
 assign add_23_2_n_26 = ~({in1[8]} & {in2[17]});
 assign add_23_2_n_25 = ({in1[8]} & {in2[27]});
 assign add_23_2_n_24 = ~({in1[3]} | {in2[3]});
 assign add_23_2_n_23 = ~({in1[3]} & {in2[3]});
 assign add_23_2_n_22 = ~({in1[8]} | {in2[23]});
 assign add_23_2_n_21 = ~({in1[8]} | {in2[16]});
 assign add_23_2_n_20 = ({in1[8]} | {in2[28]});
 assign add_23_2_n_19 = ~({in1[2]} & {in2[2]});
 assign add_23_2_n_17 = ~({in1[8]} & {in2[20]});
 assign add_23_2_n_16 = ~({in1[8]} & {in2[14]});
 assign add_23_2_n_15 = ~({in1[8]} & {in2[16]});
 assign add_23_2_n_14 = ~({in1[8]} | {in2[17]});
 assign add_23_2_n_13 = ~({in1[8]} & {in2[22]});
 assign add_23_2_n_12 = ~({in1[8]} & {in2[24]});
 assign add_23_2_n_11 = ~({in1[8]} | {in2[14]});
 assign add_23_2_n_10 = ~({in1[8]} | {in2[24]});
 assign add_23_2_n_9 = ~({in1[8]} | {in2[13]});
 assign add_23_2_n_8 = ~(n_66 & n_42);
 assign add_23_2_n_7 = ~({in1[8]} | {in2[18]});
 assign add_23_2_n_6 = ~({in1[8]} | {in2[19]});
 assign add_23_2_n_5 = ~({in1[8]} & {in2[8]});
 assign add_23_2_n_4 = ~({in1[8]} | {in2[25]});
 assign add_23_2_n_3 = ~({in1[7]} | {in2[7]});
 assign add_23_2_n_2 = ~({in1[8]} | {in2[27]});
 assign add_23_2_n_1 = ~({in1[4]} & {in2[4]});
 assign add_23_2_n_0 = ~({in1[8]} | {in2[22]});
 assign add_23_2_n_115 = ~n_115;
 assign add_23_2_n_117 = ~n_118;
 assign n_110 = ~(n_122 | (n_120 | ~add_23_2_n_16));
 assign n_111 = ~(n_121 | (n_119 | ~add_23_2_n_13));
 assign n_114 = ~(add_23_2_n_55 & add_23_2_n_12);
 assign n_115 = ~(add_23_2_n_52 & add_23_2_n_5);
 assign n_116 = (add_23_2_n_49 & add_23_2_n_39);
 assign n_117 = (add_23_2_n_28 & add_23_2_n_30);
 assign n_118 = ~(add_23_2_n_26 & add_23_2_n_15);
 assign n_119 = ~(add_23_2_n_50 & add_23_2_n_17);
 assign n_120 = ~(add_23_2_n_54 & add_23_2_n_47);
 assign n_121 = ~(add_23_2_n_53 & (add_23_2_n_117 & n_116));
 assign n_122 = ~(add_23_2_n_57 & (add_23_2_n_115 & n_117));
endmodule

