/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:10:45 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_div_cynw_cm_float_mul_ieee_E8_M23_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__46,
	inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49,
	inst_cellmath__51;
wire N440,N441,N442,N443,N444,N445,N446 
	,N447,N448,N449,N450,N461,N462,N463,N469 
	,N470,N1053,N1054,N1861,N1862,N1863,N1864;
cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I0 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw3815070899_bdw cynw_cm_float_mul_ieee_I1 (.inst_cellmath__19__2__out0(inst_cellmath__19), .inst_cellmath__19__2__in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I2 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0(inst_cellmath__19), .inst_cellmath__21_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw3815070899_bdw cynw_cm_float_mul_ieee_I3 (.inst_cellmath__13__1__out0(inst_cellmath__13), .inst_cellmath__13__1__in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw3815070899_bdw cynw_cm_float_mul_ieee_I4 (.inst_cellmath__26__9__out0({N441}), .inst_cellmath__26__9__in0(inst_cellmath__21), .inst_cellmath__26__9__in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I5 (.inst_cellmath__10_0_out0(inst_cellmath__10), .inst_cellmath__10_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw3815070899_bdw cynw_cm_float_mul_ieee_I6 (.inst_cellmath__12__0__out0(inst_cellmath__12), .inst_cellmath__12__0__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I7 (.inst_cellmath__14_0_out0(inst_cellmath__14), .inst_cellmath__14_0_in0(inst_cellmath__12), .inst_cellmath__14_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw3815070899_bdw cynw_cm_float_mul_ieee_I8 (.inst_cellmath__20__3__out0(inst_cellmath__20), .inst_cellmath__20__3__in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw3815070899_bdw cynw_cm_float_mul_ieee_I9 (.inst_cellmath__26__8__out0({N440}), .inst_cellmath__26__8__in0(inst_cellmath__20), .inst_cellmath__26__8__in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I10 (.inst_cellmath__15_0_out0(inst_cellmath__15), .inst_cellmath__15_0_in0(inst_cellmath__12), .inst_cellmath__15_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I11 (.inst_cellmath__22_0_out0(inst_cellmath__22), .inst_cellmath__22_0_in0(inst_cellmath__19), .inst_cellmath__22_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw3815070899_bdw cynw_cm_float_mul_ieee_I12 (.inst_cellmath__26_1_out0(inst_cellmath__26), .inst_cellmath__26_1_in0({N441}), .inst_cellmath__26_1_in1({N440}), .inst_cellmath__26_1_in2(inst_cellmath__22), .inst_cellmath__26_1_in3(inst_cellmath__15));
cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I13 (.inst_cellmath__23_0_out0(inst_cellmath__23), .inst_cellmath__23_0_in0(b_sign), .inst_cellmath__23_0_in1(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I14 (.inst_cellmath__41_0_out0(x[31]), .inst_cellmath__41_0_in0(inst_cellmath__26), .inst_cellmath__41_0_in1(inst_cellmath__23), .inst_cellmath__41_0_in2(inst_cellmath__22), .inst_cellmath__41_0_in3(inst_cellmath__15), .inst_cellmath__41_0_in4(b_sign), .inst_cellmath__41_0_in5(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I15 (.inst_cellmath__24_0_out0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}), .inst_cellmath__24_0_in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__24_0_in1({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I16 (.inst_cellmath__25_0_out0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24], inst_cellmath__25[23], inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}), .inst_cellmath__25_0_in0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I17 (.inst_cellmath__45_0_out0({inst_cellmath__45[24], inst_cellmath__45[23], inst_cellmath__45[22], inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__45_0_in0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw3815070899_bdw cynw_cm_float_mul_ieee_I18 (.inst_cellmath__5_1_out0(inst_cellmath__5), .inst_cellmath__5_1_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw3815070899_bdw cynw_cm_float_mul_ieee_I19 (.inst_cellmath__44__31__out0({N446}), .inst_cellmath__44__31__in0(inst_cellmath__5), .inst_cellmath__44__31__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I20 (.inst_cellmath__6_0_out0(inst_cellmath__6), .inst_cellmath__6_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw3815070899_bdw cynw_cm_float_mul_ieee_I21 (.inst_cellmath__44__30__out0({N445}), .inst_cellmath__44__30__in0(inst_cellmath__6), .inst_cellmath__44__30__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I22 (.inst_cellmath__8_0_out0(inst_cellmath__8), .inst_cellmath__8_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I23 (.inst_cellmath__4_0_out0(inst_cellmath__4), .inst_cellmath__4_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I24 (.inst_cellmath__34_0_out0(inst_cellmath__34), .inst_cellmath__34_0_in0({inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw3815070899_bdw cynw_cm_float_mul_ieee_I25 (.inst_cellmath__44__29__out0({N443}), .inst_cellmath__44__29__in0(inst_cellmath__34), .inst_cellmath__44__29__in1({inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw3815070899_bdw cynw_cm_float_mul_ieee_I26 (.inst_cellmath__44__28__out0({N444}), .inst_cellmath__44__28__in0({N443}), .inst_cellmath__44__28__in1(inst_cellmath__4));
cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw3815070899_bdw cynw_cm_float_mul_ieee_I27 (.inst_cellmath__44__27__out0({N447}), .inst_cellmath__44__27__in0(inst_cellmath__8), .inst_cellmath__44__27__in1({N446}), .inst_cellmath__44__27__in2({N445}), .inst_cellmath__44__27__in3({N444}));
cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw3815070899_bdw cynw_cm_float_mul_ieee_I28 (.inst_cellmath__44__26__out0({N448}), .inst_cellmath__44__26__in0({N447}), .inst_cellmath__44__26__in1({inst_cellmath__25[23]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw3815070899_bdw cynw_cm_float_mul_ieee_I29 (.inst_cellmath__44__33__out0({N449}), .inst_cellmath__44__33__in0({N446}), .inst_cellmath__44__33__in1({N445}));
cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw3815070899_bdw cynw_cm_float_mul_ieee_I30 (.inst_cellmath__44__32__out0({N450}), .inst_cellmath__44__32__in0({N449}), .inst_cellmath__44__32__in1(inst_cellmath__34));
cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I31 (.inst_cellmath__44_0_out0(inst_cellmath__44), .inst_cellmath__44_0_in0({N450}), .inst_cellmath__44_0_in1({N448}));
cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I32 (.inst_cellmath__46_0_out0(inst_cellmath__46), .inst_cellmath__46_0_in0({inst_cellmath__45[24]}), .inst_cellmath__46_0_in1(inst_cellmath__44));
cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I33 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__46), .inst_cellmath__38_0_in1({inst_cellmath__24[47]}));
cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I34 (.inst_cellmath__30_0_out0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}), .inst_cellmath__30_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}), .inst_cellmath__30_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I35 (.inst_cellmath__31_0_out0({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__31_0_in0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I36 (.inst_cellmath__48_0_out0({inst_cellmath__48[9], inst_cellmath__48[8], inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__48_0_in0(inst_cellmath__38), .inst_cellmath__48_0_in1({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__48_0_in2({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
INVX2 cynw_cm_float_mul_ieee_I371 (.Y(N1861), .A(inst_cellmath__48[7]));
INVX3 cynw_cm_float_mul_ieee_I372 (.Y(N1862), .A(N1861));
INVX1 cynw_cm_float_mul_ieee_I373 (.Y(N1863), .A(inst_cellmath__48[5]));
INVX2 cynw_cm_float_mul_ieee_I374 (.Y(N1864), .A(N1863));
INVXL cynw_cm_float_mul_ieee_I136 (.Y(N1053), .A(inst_cellmath__48[2]));
INVX2 cynw_cm_float_mul_ieee_I137 (.Y(N1054), .A(N1053));
cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw3815070899_bdw cynw_cm_float_mul_ieee_I37 (.inst_cellmath__51__49__out0({N461}), .inst_cellmath__51__49__in0({inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], N1054, inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw3815070899_bdw cynw_cm_float_mul_ieee_I38 (.inst_cellmath__51__48__out0({N462}), .inst_cellmath__51__48__in0({N461}), .inst_cellmath__51__48__in1({inst_cellmath__48[8]}));
cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I39 (.inst_cellmath__51_0_out0(inst_cellmath__51), .inst_cellmath__51_0_in0({N462}), .inst_cellmath__51_0_in1({inst_cellmath__48[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I40 (.inst_cellmath__28_0_out0(inst_cellmath__28), .inst_cellmath__28_0_in0(inst_cellmath__20), .inst_cellmath__28_0_in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I41 (.inst_cellmath__27_0_out0(inst_cellmath__27), .inst_cellmath__27_0_in0(inst_cellmath__21), .inst_cellmath__27_0_in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw3815070899_bdw cynw_cm_float_mul_ieee_I42 (.inst_cellmath__50__50__out0({N463}), .inst_cellmath__50__50__in0({inst_cellmath__48[9], inst_cellmath__48[8], N1862, inst_cellmath__48[6], N1864, inst_cellmath__48[4], inst_cellmath__48[3], N1054, inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw3815070899_bdw cynw_cm_float_mul_ieee_I43 (.inst_cellmath__49_1_out0(inst_cellmath__49), .inst_cellmath__49_1_in0(inst_cellmath__51), .inst_cellmath__49_1_in1({N463}), .inst_cellmath__49_1_in2({inst_cellmath__48[9]}), .inst_cellmath__49_1_in3(inst_cellmath__28), .inst_cellmath__49_1_in4(inst_cellmath__27), .inst_cellmath__49_1_in5(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw3815070899_bdw cynw_cm_float_mul_ieee_I44 (.inst_cellmath__37__43__out0({N470}), .inst_cellmath__37__43__in0(inst_cellmath__27), .inst_cellmath__37__43__in1(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw3815070899_bdw cynw_cm_float_mul_ieee_I45 (.inst_cellmath__32__11__out0({N442}), .inst_cellmath__32__11__in0({inst_cellmath__30[8], inst_cellmath__30[7]}));
cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw3815070899_bdw cynw_cm_float_mul_ieee_I46 (.inst_cellmath__32__10__out0(inst_cellmath__32), .inst_cellmath__32__10__in0({N442}), .inst_cellmath__32__10__in1({inst_cellmath__30[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw3815070899_bdw cynw_cm_float_mul_ieee_I47 (.inst_cellmath__37__42__out0({N469}), .inst_cellmath__37__42__in0(inst_cellmath__32), .inst_cellmath__37__42__in1(inst_cellmath__28));
cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I48 (.inst_cellmath__7_0_out0(inst_cellmath__7), .inst_cellmath__7_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I49 (.inst_cellmath__42_0_out0(inst_cellmath__42), .inst_cellmath__42_0_in0(inst_cellmath__7), .inst_cellmath__42_0_in1(inst_cellmath__6), .inst_cellmath__42_0_in2(inst_cellmath__5), .inst_cellmath__42_0_in3(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I50 (.inst_cellmath__52_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__52_0_in0(inst_cellmath__49), .inst_cellmath__52_0_in1({N1862, inst_cellmath__48[6], N1864, inst_cellmath__48[4], inst_cellmath__48[3], N1054, inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__52_0_in2(inst_cellmath__42), .inst_cellmath__52_0_in3({N470}), .inst_cellmath__52_0_in4({N469}));
cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw3815070899_bdw cynw_cm_float_mul_ieee_I51 (.inst_cellmath__47_0_out0(inst_cellmath__47), .inst_cellmath__47_0_in0(inst_cellmath__42), .inst_cellmath__47_0_in1(inst_cellmath__32), .inst_cellmath__47_0_in2(inst_cellmath__28), .inst_cellmath__47_0_in3(inst_cellmath__27), .inst_cellmath__47_0_in4(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw3815070899_bdw cynw_cm_float_mul_ieee_I52 (.inst_cellmath__53_U_out0({x[22]}), .inst_cellmath__53_U_in0(inst_cellmath__49), .inst_cellmath__53_U_in1(inst_cellmath__47), .inst_cellmath__53_U_in2({inst_cellmath__45[22]}), .inst_cellmath__53_U_in3(inst_cellmath__44), .inst_cellmath__53_U_in4(inst_cellmath__26), .inst_cellmath__53_U_in5({inst_cellmath__25[46]}));
cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw3815070899_bdw cynw_cm_float_mul_ieee_I53 (.inst_cellmath__53_M_out0({x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__53_M_in0(inst_cellmath__49), .inst_cellmath__53_M_in1(inst_cellmath__47), .inst_cellmath__53_M_in2({inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__53_M_in3(inst_cellmath__44), .inst_cellmath__53_M_in4(inst_cellmath__26), .inst_cellmath__53_M_in5({inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}), .inst_cellmath__53_M_in6(inst_cellmath__22), .inst_cellmath__53_M_in7(inst_cellmath__15), .inst_cellmath__53_M_in8({b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__53_M_in9({a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw3815070899_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2X1 inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[0]), .B(inst_cellmath__17_0_in0[1]));
NAND2XL inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[6]));
NAND2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[5]), .B(inst_cellmath__17_0_in0[4]));
NAND2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[3]), .B(inst_cellmath__17_0_in0[2]));
NOR2XL inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw3815070899_bdw (
	inst_cellmath__19__2__out0,
	inst_cellmath__19__2__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19__2__out0;
input [22:0] inst_cellmath__19__2__in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48;
NOR2XL inst_cellmath__19__2__I0 (.Y(N26), .A(inst_cellmath__19__2__in0[0]), .B(inst_cellmath__19__2__in0[1]));
NOR2XL inst_cellmath__19__2__I1 (.Y(N27), .A(inst_cellmath__19__2__in0[22]), .B(inst_cellmath__19__2__in0[21]));
NOR2XL inst_cellmath__19__2__I2 (.Y(N28), .A(inst_cellmath__19__2__in0[20]), .B(inst_cellmath__19__2__in0[19]));
NOR2XL inst_cellmath__19__2__I3 (.Y(N29), .A(inst_cellmath__19__2__in0[18]), .B(inst_cellmath__19__2__in0[17]));
NOR2XL inst_cellmath__19__2__I4 (.Y(N30), .A(inst_cellmath__19__2__in0[16]), .B(inst_cellmath__19__2__in0[15]));
NOR2XL inst_cellmath__19__2__I5 (.Y(N31), .A(inst_cellmath__19__2__in0[14]), .B(inst_cellmath__19__2__in0[13]));
NOR2XL inst_cellmath__19__2__I6 (.Y(N32), .A(inst_cellmath__19__2__in0[12]), .B(inst_cellmath__19__2__in0[11]));
NOR2XL inst_cellmath__19__2__I7 (.Y(N33), .A(inst_cellmath__19__2__in0[10]), .B(inst_cellmath__19__2__in0[9]));
NOR2XL inst_cellmath__19__2__I8 (.Y(N34), .A(inst_cellmath__19__2__in0[8]), .B(inst_cellmath__19__2__in0[7]));
NOR2XL inst_cellmath__19__2__I9 (.Y(N35), .A(inst_cellmath__19__2__in0[6]), .B(inst_cellmath__19__2__in0[5]));
NOR2XL inst_cellmath__19__2__I10 (.Y(N36), .A(inst_cellmath__19__2__in0[4]), .B(inst_cellmath__19__2__in0[3]));
INVXL inst_cellmath__19__2__I11 (.Y(N37), .A(inst_cellmath__19__2__in0[2]));
NAND2XL inst_cellmath__19__2__I12 (.Y(N38), .A(N37), .B(N26));
NAND2XL inst_cellmath__19__2__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__19__2__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__19__2__I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__19__2__I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__19__2__I17 (.Y(N43), .A(N35), .B(N36));
NOR2XL inst_cellmath__19__2__I18 (.Y(N44), .A(N38), .B(N39));
NOR2XL inst_cellmath__19__2__I19 (.Y(N45), .A(N40), .B(N41));
NAND2XL inst_cellmath__19__2__I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__19__2__I169 (.Y(N48), .A(N42), .B(N43));
NOR2XL inst_cellmath__19__2__I23 (.Y(inst_cellmath__19__2__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw3815070899_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input  inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1;
AND2XL inst_cellmath__21_0_I0 (.Y(inst_cellmath__21_0_out0), .A(inst_cellmath__21_0_in1), .B(inst_cellmath__21_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw3815070899_bdw (
	inst_cellmath__13__1__out0,
	inst_cellmath__13__1__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__13__1__out0;
input [7:0] inst_cellmath__13__1__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2X1 inst_cellmath__13__1__I0 (.Y(N11), .A(inst_cellmath__13__1__in0[0]), .B(inst_cellmath__13__1__in0[1]));
NOR2X1 inst_cellmath__13__1__I1 (.Y(N12), .A(inst_cellmath__13__1__in0[7]), .B(inst_cellmath__13__1__in0[6]));
NOR2XL inst_cellmath__13__1__I2 (.Y(N13), .A(inst_cellmath__13__1__in0[5]), .B(inst_cellmath__13__1__in0[4]));
NOR2XL inst_cellmath__13__1__I3 (.Y(N14), .A(inst_cellmath__13__1__in0[3]), .B(inst_cellmath__13__1__in0[2]));
NAND2X1 inst_cellmath__13__1__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__13__1__I5 (.Y(N16), .A(N13), .B(N14));
NOR2X1 inst_cellmath__13__1__I6 (.Y(inst_cellmath__13__1__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw3815070899_bdw (
	inst_cellmath__26__9__out0,
	inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__9__out0;
input  inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1;
wire N19;
NAND2X2 inst_cellmath__26__9__I4 (.Y(N19), .A(inst_cellmath__26__9__in1), .B(inst_cellmath__26__9__in0));
INVXL inst_cellmath__26__9__I5 (.Y(inst_cellmath__26__9__out0[0]), .A(N19));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw3815070899_bdw (
	inst_cellmath__10_0_out0,
	inst_cellmath__10_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__10_0_out0;
input [7:0] inst_cellmath__10_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2X1 inst_cellmath__10_0_I0 (.Y(N11), .A(inst_cellmath__10_0_in0[0]), .B(inst_cellmath__10_0_in0[1]));
NAND2XL inst_cellmath__10_0_I1 (.Y(N12), .A(inst_cellmath__10_0_in0[7]), .B(inst_cellmath__10_0_in0[6]));
NAND2XL inst_cellmath__10_0_I2 (.Y(N13), .A(inst_cellmath__10_0_in0[5]), .B(inst_cellmath__10_0_in0[4]));
NAND2XL inst_cellmath__10_0_I3 (.Y(N14), .A(inst_cellmath__10_0_in0[3]), .B(inst_cellmath__10_0_in0[2]));
NOR2XL inst_cellmath__10_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__10_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__10_0_I6 (.Y(inst_cellmath__10_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw3815070899_bdw (
	inst_cellmath__12__0__out0,
	inst_cellmath__12__0__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__12__0__out0;
input [22:0] inst_cellmath__12__0__in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48;
NOR2XL inst_cellmath__12__0__I0 (.Y(N26), .A(inst_cellmath__12__0__in0[0]), .B(inst_cellmath__12__0__in0[1]));
NOR2XL inst_cellmath__12__0__I1 (.Y(N27), .A(inst_cellmath__12__0__in0[22]), .B(inst_cellmath__12__0__in0[21]));
NOR2XL inst_cellmath__12__0__I2 (.Y(N28), .A(inst_cellmath__12__0__in0[20]), .B(inst_cellmath__12__0__in0[19]));
NOR2XL inst_cellmath__12__0__I3 (.Y(N29), .A(inst_cellmath__12__0__in0[18]), .B(inst_cellmath__12__0__in0[17]));
NOR2XL inst_cellmath__12__0__I4 (.Y(N30), .A(inst_cellmath__12__0__in0[16]), .B(inst_cellmath__12__0__in0[15]));
NOR2XL inst_cellmath__12__0__I5 (.Y(N31), .A(inst_cellmath__12__0__in0[14]), .B(inst_cellmath__12__0__in0[13]));
NOR2XL inst_cellmath__12__0__I6 (.Y(N32), .A(inst_cellmath__12__0__in0[12]), .B(inst_cellmath__12__0__in0[11]));
NOR2XL inst_cellmath__12__0__I7 (.Y(N33), .A(inst_cellmath__12__0__in0[10]), .B(inst_cellmath__12__0__in0[9]));
NOR2XL inst_cellmath__12__0__I8 (.Y(N34), .A(inst_cellmath__12__0__in0[8]), .B(inst_cellmath__12__0__in0[7]));
NOR2XL inst_cellmath__12__0__I9 (.Y(N35), .A(inst_cellmath__12__0__in0[6]), .B(inst_cellmath__12__0__in0[5]));
NOR2XL inst_cellmath__12__0__I10 (.Y(N36), .A(inst_cellmath__12__0__in0[4]), .B(inst_cellmath__12__0__in0[3]));
INVXL inst_cellmath__12__0__I11 (.Y(N37), .A(inst_cellmath__12__0__in0[2]));
NAND2XL inst_cellmath__12__0__I12 (.Y(N38), .A(N37), .B(N26));
NAND2XL inst_cellmath__12__0__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__12__0__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__12__0__I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__12__0__I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__12__0__I17 (.Y(N43), .A(N35), .B(N36));
NOR2XL inst_cellmath__12__0__I18 (.Y(N44), .A(N38), .B(N39));
NOR2XL inst_cellmath__12__0__I19 (.Y(N45), .A(N40), .B(N41));
NAND2XL inst_cellmath__12__0__I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__12__0__I169 (.Y(N48), .A(N42), .B(N43));
NOR2XL inst_cellmath__12__0__I23 (.Y(inst_cellmath__12__0__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw3815070899_bdw (
	inst_cellmath__14_0_out0,
	inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__14_0_out0;
input  inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1;
AND2XL inst_cellmath__14_0_I0 (.Y(inst_cellmath__14_0_out0), .A(inst_cellmath__14_0_in1), .B(inst_cellmath__14_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw3815070899_bdw (
	inst_cellmath__20__3__out0,
	inst_cellmath__20__3__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__20__3__out0;
input [7:0] inst_cellmath__20__3__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2X1 inst_cellmath__20__3__I0 (.Y(N11), .A(inst_cellmath__20__3__in0[0]), .B(inst_cellmath__20__3__in0[1]));
NOR2X1 inst_cellmath__20__3__I1 (.Y(N12), .A(inst_cellmath__20__3__in0[7]), .B(inst_cellmath__20__3__in0[6]));
NOR2XL inst_cellmath__20__3__I2 (.Y(N13), .A(inst_cellmath__20__3__in0[5]), .B(inst_cellmath__20__3__in0[4]));
NOR2XL inst_cellmath__20__3__I3 (.Y(N14), .A(inst_cellmath__20__3__in0[3]), .B(inst_cellmath__20__3__in0[2]));
NAND2X1 inst_cellmath__20__3__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__20__3__I5 (.Y(N16), .A(N13), .B(N14));
NOR2X1 inst_cellmath__20__3__I6 (.Y(inst_cellmath__20__3__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw3815070899_bdw (
	inst_cellmath__26__8__out0,
	inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__8__out0;
input  inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1;
AND2XL inst_cellmath__26__8__I0 (.Y(inst_cellmath__26__8__out0[0]), .A(inst_cellmath__26__8__in0), .B(inst_cellmath__26__8__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw3815070899_bdw (
	inst_cellmath__15_0_out0,
	inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__15_0_out0;
input  inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1;
wire N5;
INVXL inst_cellmath__15_0_I0 (.Y(N5), .A(inst_cellmath__15_0_in1));
NOR2X2 inst_cellmath__15_0_I1 (.Y(inst_cellmath__15_0_out0), .A(N5), .B(inst_cellmath__15_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw3815070899_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__22_0_out0;
input  inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1;
wire N5;
INVXL inst_cellmath__22_0_I0 (.Y(N5), .A(inst_cellmath__22_0_in1));
NOR2X2 inst_cellmath__22_0_I1 (.Y(inst_cellmath__22_0_out0), .A(N5), .B(inst_cellmath__22_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw3815070899_bdw (
	inst_cellmath__26_1_out0,
	inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1,
	inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__26_1_out0;
input [0:0] inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1;
input  inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3;
wire N7,N8,N9,N10;
NOR2XL inst_cellmath__26_1_I0 (.Y(N7), .A(inst_cellmath__26_1_in3), .B(inst_cellmath__26_1_in2));
INVXL inst_cellmath__26_1_I1 (.Y(N8), .A(N7));
NOR2XL inst_cellmath__26_1_I2 (.Y(N9), .A(N8), .B(inst_cellmath__26_1_in0[0]));
INVXL inst_cellmath__26_1_I3 (.Y(N10), .A(inst_cellmath__26_1_in1[0]));
NAND2XL inst_cellmath__26_1_I4 (.Y(inst_cellmath__26_1_out0), .A(N10), .B(N9));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw3815070899_bdw (
	inst_cellmath__23_0_out0,
	inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__23_0_out0;
input  inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1;
wire N2,N6;
INVXL inst_cellmath__23_0_I1 (.Y(N6), .A(inst_cellmath__23_0_in1));
MXI2XL inst_cellmath__23_0_I2 (.Y(N2), .A(N6), .B(inst_cellmath__23_0_in1), .S0(inst_cellmath__23_0_in0));
btree_10_bdw3815070899_bdw inst_cellmath__23_0_I3 (.Y(inst_cellmath__23_0_out0), .A(N2));
endmodule

`ifdef btree_10_bdw3815070899_bdw_COMPILED
`else
`define btree_10_bdw3815070899_bdw_COMPILED
module btree_10_bdw3815070899_bdw (
	A,
	Y
	); /* architecture "gate_level" */ 
input  A;
output  Y;
assign Y = A;
endmodule
`endif //  `ifdef btree_10_bdw3815070899_bdw_COMPILED

module cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw3815070899_bdw (
	inst_cellmath__41_0_out0,
	inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__41_0_out0;
input  inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5;
wire N15,N18,N19;
NAND2BXL inst_cellmath__41_0_I12 (.Y(N15), .AN(inst_cellmath__41_0_in4), .B(inst_cellmath__41_0_in2));
MXI2XL inst_cellmath__41_0_I13 (.Y(N18), .A(N15), .B(inst_cellmath__41_0_in5), .S0(inst_cellmath__41_0_in3));
INVXL inst_cellmath__41_0_I6 (.Y(N19), .A(inst_cellmath__41_0_in1));
MXI2XL inst_cellmath__41_0_I11 (.Y(inst_cellmath__41_0_out0), .A(N19), .B(N18), .S0(inst_cellmath__41_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw3815070899_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1;
wire N383,N385,N387,N389,N391,N393,N395 
	,N397,N399,N401,N403,N405,N407,N409,N411 
	,N413,N415,N417,N419,N421,N423,N425,N427 
	,N440,N442,N444,N446,N448,N450,N452,N454 
	,N456,N458,N460,N462,N464,N466,N468,N470 
	,N472,N474,N476,N478,N480,N482,N484,N486 
	,N499,N501,N503,N505,N507,N509,N511,N513 
	,N515,N517,N519,N521,N523,N525,N527,N529 
	,N531,N533,N535,N537,N539,N541,N543,N545 
	,N558,N560,N562,N564,N566,N568,N570,N572 
	,N574,N576,N578,N580,N582,N584,N586,N588 
	,N590,N592,N594,N596,N598,N600,N602,N604 
	,N617,N619,N621,N623,N625,N627,N629,N631 
	,N633,N635,N637,N639,N641,N643,N645,N647 
	,N649,N651,N653,N655,N657,N659,N661,N663 
	,N676,N678,N680,N682,N684,N686,N688,N690 
	,N692,N694,N696,N698,N700,N702,N704,N706 
	,N708,N710,N712,N714,N716,N718,N720,N722 
	,N735,N737,N739,N741,N743,N745,N747,N749 
	,N751,N753,N755,N757,N759,N761,N763,N765 
	,N767,N769,N771,N773,N775,N777,N779,N781 
	,N794,N796,N798,N800,N802,N804,N806,N808 
	,N810,N812,N814,N816,N818,N820,N822,N824 
	,N826,N828,N830,N832,N834,N836,N838,N840 
	,N853,N855,N857,N859,N861,N863,N865,N867 
	,N869,N871,N873,N875,N877,N879,N881,N883 
	,N885,N887,N889,N891,N893,N895,N897,N899 
	,N912,N914,N916,N918,N920,N922,N924,N926 
	,N928,N930,N932,N934,N936,N938,N940,N942 
	,N944,N946,N948,N950,N952,N954,N956,N958 
	,N971,N973,N975,N977,N979,N981,N983,N985 
	,N987,N989,N991,N993,N995,N997,N999,N1001 
	,N1003,N1005,N1007,N1009,N1011,N1013,N1015,N1017 
	,N1030,N1032,N1034,N1036,N1038,N1040,N1042,N1044 
	,N1046,N1048,N1050,N1052,N1054,N1056,N1058,N1060 
	,N1062,N1064,N1066,N1068,N1070,N1072,N1074,N1076 
	,N1089,N1091,N1093,N1095,N1097,N1099,N1101,N1103 
	,N1105,N1107,N1109,N1111,N1113,N1115,N1117,N1119 
	,N1121,N1123,N1125,N1127,N1129,N1131,N1133,N1135 
	,N1148,N1150,N1152,N1154,N1156,N1158,N1160,N1162 
	,N1164,N1166,N1168,N1170,N1172,N1174,N1176,N1178 
	,N1180,N1182,N1184,N1186,N1188,N1190,N1192,N1194 
	,N1207,N1209,N1211,N1213,N1215,N1217,N1219,N1221 
	,N1223,N1225,N1227,N1229,N1231,N1233,N1235,N1237 
	,N1239,N1241,N1243,N1245,N1247,N1249,N1251,N1253 
	,N1266,N1268,N1270,N1272,N1274,N1276,N1278,N1280 
	,N1282,N1284,N1286,N1288,N1290,N1292,N1294,N1296 
	,N1298,N1300,N1302,N1304,N1306,N1308,N1310,N1312 
	,N1325,N1327,N1329,N1331,N1333,N1335,N1337,N1339 
	,N1341,N1343,N1345,N1347,N1349,N1351,N1353,N1355 
	,N1357,N1359,N1361,N1363,N1365,N1367,N1369,N1371 
	,N1384,N1386,N1388,N1390,N1392,N1394,N1396,N1398 
	,N1400,N1402,N1404,N1406,N1408,N1410,N1412,N1414 
	,N1416,N1418,N1420,N1422,N1424,N1426,N1428,N1430 
	,N1443,N1445,N1447,N1449,N1451,N1453,N1455,N1457 
	,N1459,N1461,N1463,N1465,N1467,N1469,N1471,N1473 
	,N1475,N1477,N1479,N1481,N1483,N1485,N1487,N1489 
	,N1502,N1504,N1506,N1508,N1510,N1512,N1514,N1516 
	,N1518,N1520,N1522,N1524,N1526,N1528,N1530,N1532 
	,N1534,N1536,N1538,N1540,N1542,N1544,N1546,N1548 
	,N1561,N1563,N1565,N1567,N1569,N1571,N1573,N1575 
	,N1577,N1579,N1581,N1583,N1585,N1587,N1589,N1591 
	,N1593,N1595,N1597,N1599,N1601,N1603,N1605,N1607 
	,N1620,N1622,N1624,N1626,N1628,N1630,N1632,N1634 
	,N1636,N1638,N1640,N1642,N1644,N1646,N1648,N1650 
	,N1652,N1654,N1656,N1658,N1660,N1662,N1664,N1666 
	,N1679,N1681,N1683,N1685,N1687,N1689,N1691,N1693 
	,N1695,N1697,N1699,N1701,N1703,N1705,N1707,N1709 
	,N1711,N1713,N1715,N1717,N1719,N1721,N1723,N1725 
	,N1734,N1736,N1738,N1740,N1742,N1744,N1746,N1748 
	,N1750,N1752,N1754,N1756,N1758,N1760,N1762,N1764 
	,N1766,N1768,N1770,N1772,N1774,N1776,N1778,N1782 
	,N1783,N1784,N1785,N1786,N1787,N1788,N1789,N1790 
	,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798 
	,N1799,N1800,N1801,N1802,N1803,N1804,N1805,N1806 
	,N1807,N1808,N1809,N1810,N1811,N1812,N1813,N1814 
	,N1815,N1816,N1817,N1818,N1819,N1820,N1821,N1822 
	,N1823,N1824,N1825,N1826,N1827,N1828,N1829,N1830 
	,N1831,N1832,N1833,N1834,N1835,N1836,N1837,N1838 
	,N1839,N1840,N1841,N1842,N1843,N1844,N1845,N1846 
	,N1847,N1848,N1849,N1850,N1851,N1852,N1853,N1854 
	,N1855,N1856,N1857,N1858,N1859,N1860,N1861,N1862 
	,N1863,N1864,N1865,N1866,N1867,N1868,N1869,N1870 
	,N1871,N1872,N1873,N1874,N1875,N1876,N1877,N1878 
	,N1879,N1880,N1881,N1882,N1883,N1884,N1885,N1886 
	,N1887,N1888,N1889,N1890,N1891,N1892,N1893,N1894 
	,N1895,N1896,N1897,N1898,N1899,N1900,N1901,N1902 
	,N1903,N1904,N1905,N1906,N1907,N1908,N1909,N1910 
	,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918 
	,N1919,N1920,N1921,N1922,N1923,N1924,N1925,N1926 
	,N1927,N1928,N1929,N1930,N1931,N1932,N1933,N1934 
	,N1935,N1936,N1937,N1938,N1939,N1940,N1941,N1942 
	,N1943,N1944,N1945,N1946,N1947,N1948,N1949,N1950 
	,N1951,N1952,N1953,N1954,N1955,N1956,N1957,N1958 
	,N1959,N1960,N1961,N1962,N1963,N1964,N1965,N1966 
	,N1967,N1968,N1969,N1970,N1971,N1972,N1973,N1974 
	,N1975,N1976,N1977,N1978,N1979,N1980,N1981,N1982 
	,N1983,N1984,N1985,N1986,N1987,N1988,N1989,N1990 
	,N1991,N1992,N1993,N1994,N1995,N1996,N1997,N1998 
	,N1999,N2000,N2001,N2002,N2003,N2004,N2005,N2006 
	,N2007,N2008,N2009,N2010,N2011,N2012,N2013,N2014 
	,N2015,N2016,N2017,N2018,N2019,N2020,N2021,N2022 
	,N2023,N2024,N2025,N2026,N2027,N2028,N2029,N2030 
	,N2031,N2032,N2033,N2034,N2035,N2036,N2037,N2038 
	,N2039,N2040,N2041,N2042,N2043,N2044,N2045,N2046 
	,N2047,N2048,N2049,N2050,N2051,N2052,N2053,N2054 
	,N2055,N2056,N2057,N2058,N2059,N2060,N2061,N2062 
	,N2063,N2064,N2065,N2066,N2067,N2068,N2069,N2070 
	,N2071,N2072,N2073,N2074,N2075,N2076,N2077,N2078 
	,N2079,N2080,N2081,N2082,N2083,N2084,N2085,N2086 
	,N2087,N2088,N2089,N2090,N2091,N2092,N2093,N2094 
	,N2095,N2096,N2097,N2098,N2099,N2100,N2101,N2102 
	,N2103,N2104,N2105,N2106,N2107,N2108,N2109,N2110 
	,N2111,N2112,N2113,N2114,N2115,N2116,N2117,N2118 
	,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126 
	,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134 
	,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142 
	,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150 
	,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158 
	,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166 
	,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174 
	,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182 
	,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190 
	,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198 
	,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206 
	,N2207,N2208,N2209,N2210,N2211,N2212,N2213,N2214 
	,N2215,N2216,N2217,N2218,N2219,N2220,N2221,N2222 
	,N2223,N2224,N2225,N2226,N2227,N2228,N2229,N2230 
	,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238 
	,N2239,N2240,N2241,N2242,N2243,N2244,N2245,N2246 
	,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254 
	,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262 
	,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270 
	,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278 
	,N2279,N2280,N2281,N2282,N2283,N2284,N2285,N2286 
	,N2287,N2288,N2289,N2290,N2291,N2292,N2293,N2294 
	,N2295,N2296,N2297,N2298,N2299,N2300,N2301,N2302 
	,N2303,N2304,N2305,N2306,N2307,N2308,N2309,N2310 
	,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318 
	,N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326 
	,N2327,N2328,N2329,N2330,N2331,N2332,N2333,N2334 
	,N2335,N2336,N2337,N2338,N2339,N2340,N2341,N2342 
	,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350 
	,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358 
	,N2359,N2360,N2361,N2362,N2363,N2364,N2365,N2366 
	,N2367,N2368,N2369,N2370,N2371,N2372,N2373,N2374 
	,N2375,N2376,N2377,N2378,N2379,N2380,N2381,N2382 
	,N2383,N2384,N2385,N2386,N2387,N2388,N2389,N2390 
	,N2391,N2392,N2393,N2394,N2395,N2396,N2397,N2398 
	,N2399,N2400,N2401,N2402,N2403,N2404,N2405,N2406 
	,N2407,N2408,N2409,N2410,N2411,N2412,N2413,N2414 
	,N2415,N2416,N2417,N2418,N2419,N2420,N2421,N2422 
	,N2423,N2424,N2425,N2426,N2427,N2428,N2429,N2430 
	,N2431,N2432,N2433,N2434,N2435,N2436,N2437,N2438 
	,N2439,N2440,N2441,N2442,N2443,N2444,N2445,N2446 
	,N2447,N2448,N2449,N2450,N2451,N2452,N2453,N2454 
	,N2455,N2456,N2457,N2458,N2459,N2460,N2461,N2462 
	,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470 
	,N2471,N2472,N2473,N2474,N2475,N2476,N2477,N2478 
	,N2479,N2480,N2481,N2482,N2483,N2484,N2485,N2486 
	,N2487,N2488,N2489,N2490,N2491,N2492,N2493,N2494 
	,N2495,N2496,N2497,N2498,N2499,N2500,N2501,N2502 
	,N2503,N2504,N2505,N2506,N2507,N2508,N2509,N2510 
	,N2511,N2512,N2513,N2514,N2515,N2516,N2517,N2518 
	,N2519,N2520,N2521,N2522,N2523,N2524,N2525,N2526 
	,N2527,N2528,N2529,N2530,N2531,N2532,N2533,N2534 
	,N2535,N2536,N2537,N2538,N2539,N2540,N2541,N2542 
	,N2543,N2544,N2545,N2546,N2547,N2548,N2549,N2550 
	,N2551,N2552,N2553,N2554,N2555,N2556,N2557,N2558 
	,N2559,N2560,N2561,N2562,N2563,N2564,N2565,N2566 
	,N2567,N2568,N2569,N2570,N2571,N2572,N2573,N2574 
	,N2575,N2576,N2577,N2578,N2579,N2580,N2581,N2582 
	,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590 
	,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598 
	,N2599,N2600,N2601,N2602,N2603,N2604,N2605,N2606 
	,N2607,N2608,N2609,N2610,N2611,N2612,N2613,N2614 
	,N2615,N2616,N2617,N2618,N2619,N2620,N2621,N2622 
	,N2623,N2624,N2625,N2626,N2627,N2628,N2629,N2630 
	,N2631,N2632,N2633,N2634,N2635,N2636,N2637,N2638 
	,N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646 
	,N2647,N2648,N2649,N2650,N2651,N2652,N2653,N2654 
	,N2655,N2656,N2657,N2658,N2659,N2660,N2661,N2662 
	,N2663,N2664,N2665,N2666,N2667,N2668,N2669,N2670 
	,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678 
	,N2679,N2680,N2681,N2682,N2683,N2684,N2685,N2686 
	,N2687,N2688,N2689,N2690,N2691,N2692,N2693,N2694 
	,N2695,N2696,N2697,N2698,N2699,N2700,N2701,N2702 
	,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710 
	,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718 
	,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726 
	,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734 
	,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742 
	,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750 
	,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758 
	,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2766 
	,N2767,N2768,N2769,N2770,N2771,N2772,N2773,N2774 
	,N2775,N2776,N2777,N2778,N2779,N2780,N2781,N2782 
	,N2783,N2784,N2785,N2786,N2787,N2788,N2789,N2790 
	,N2791,N2792,N2794,N2795,N2796,N2797,N2798,N2799 
	,N2800,N2801,N2802,N2803,N2804,N2805,N2806,N2807 
	,N2808,N2809,N2810,N2811,N2812,N2813,N2814,N2815 
	,N2816,N2817,N2818,N2819,N2820,N2823,N2831,N2839 
	,N2851,N2863,N2879,N2903,N2905,N2909,N2910,N2931 
	,N2955,N2959,N2960,N2985,N2994,N2997,N3000,N3003 
	,N3006,N3009,N3012,N3015,N3018,N3021,N3024,N3027 
	,N3030,N3046,N3048,N3049,N3050,N3051,N3052,N3053 
	,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061 
	,N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069 
	,N3070,N3071,N3072,N3073,N3074,N3075,N3076,N3077 
	,N3078,N3079,N3080,N3081,N3082,N3083,N3084,N3085 
	,N3086,N3087,N3088,N3089,N3090,N3091,N3092,N3093 
	,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101 
	,N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109 
	,N3110,N3113,N3117,N3118,N3121,N3122,N3127,N3129 
	,N3130,N3133,N3137,N3138,N3141,N3145,N3146,N3149 
	,N3153,N3157,N3158,N3161,N3162,N3167,N3169,N3170 
	,N3173,N3174,N3177,N3178,N3183,N3185,N3186,N3189 
	,N3190,N3193,N3194,N3199,N3205,N3206,N3215,N3246 
	,N3250,N3251,N3258,N3262,N3263,N3266,N3267,N3272 
	,N3273,N3274,N3275,N3284,N3286,N3288,N3290,N3294 
	,N3295,N3302,N3326,N3328,N3330,N3337,N3340,N3343 
	,N3346,N3349,N3352,N3355,N3358,N3361,N3364,N3367 
	,N3370,N3373,N3376,N3379,N3382,N3385,N3388,N3391 
	,N3394,N3397,N3400,N3403,N3406,N3409,N3412,N3415 
	,N3418,N3421,N3424,N3427,N3445,N3446,N3448,N3449 
	,N3451,N3452,N3454,N3455,N3457,N3458,N3460,N3461 
	,N3463,N3464,N3466,N3467,N3469,N3470,N3472,N3473 
	,N3475,N3476,N3478,N3479,N3481,N3482,N3484,N3485 
	,N3487,N3488,N3490,N3491,N3493,N3494,N3496,N3497 
	,N3499,N3500,N3502,N3503,N3505,N3623,N3632,N3690 
	,N3699,N3715,N3724,N3740,N3749,N3765,N3793,N3797 
	,N3805,N3813,N3820,N3821,N3826,N3829,N3834,N3837 
	,N3845,N3853,N3861,N3869,N3877,N3885,N3891,N3893 
	,N3900,N3901,N3909,N3917,N3925,N3933,N3941,N3949 
	,N3957,N3965,N3973,N3977,N3981,N3989,N3994,N3997 
	,N4003,N4004,N4007,N4010,N4011,N4016,N4017,N4018 
	,N4023,N4025,N4031,N4033,N4039,N4041,N4047,N4048 
	,N4053,N4055,N4063,N4068,N4070,N4071,N4078,N4079 
	,N4087,N4094,N4101,N4109,N4116,N4117,N4125,N4133 
	,N4141,N4149,N4152,N4153,N4159,N4160,N4170,N4171 
	,N4182,N4183,N4213,N4217,N4218,N4224,N4225,N4228 
	,N4244,N4245,N4248,N4252,N4253,N4256,N4260,N4261 
	,N4264,N4272,N4274,N4277,N4278,N4281,N4282,N4285 
	,N4286,N4289,N4290,N4293,N4294,N4297,N4298,N4299 
	,N4303,N4314,N4315,N4318,N4319,N4322,N4323,N4325 
	,N4328,N4329,N4334,N4335,N4338,N4339,N4344,N4346 
	,N4374,N4381,N4388,N4395,N4407,N8767;
INVX1 inst_cellmath__24_0_I2067 (.Y(N3797), .A(inst_cellmath__24_0_in1[0]));
INVXL inst_cellmath__24_0_I2063 (.Y(N3793), .A(inst_cellmath__24_0_in1[0]));
INVX2 inst_cellmath__24_0_I2075 (.Y(N3805), .A(inst_cellmath__24_0_in1[1]));
INVX2 inst_cellmath__24_0_I2083 (.Y(N3813), .A(inst_cellmath__24_0_in1[2]));
INVXL inst_cellmath__24_0_I2091 (.Y(N3821), .A(inst_cellmath__24_0_in1[3]));
INVX2 inst_cellmath__24_0_I2090 (.Y(N3820), .A(inst_cellmath__24_0_in1[3]));
INVX1 inst_cellmath__24_0_I2099 (.Y(N3829), .A(inst_cellmath__24_0_in1[4]));
INVX1 inst_cellmath__24_0_I2096 (.Y(N3826), .A(inst_cellmath__24_0_in1[4]));
INVX1 inst_cellmath__24_0_I2107 (.Y(N3837), .A(inst_cellmath__24_0_in1[5]));
INVX2 inst_cellmath__24_0_I2104 (.Y(N3834), .A(inst_cellmath__24_0_in1[5]));
INVX3 inst_cellmath__24_0_I2115 (.Y(N3845), .A(inst_cellmath__24_0_in1[6]));
INVX3 inst_cellmath__24_0_I2123 (.Y(N3853), .A(inst_cellmath__24_0_in1[7]));
INVX2 inst_cellmath__24_0_I2131 (.Y(N3861), .A(inst_cellmath__24_0_in1[8]));
INVX3 inst_cellmath__24_0_I2139 (.Y(N3869), .A(inst_cellmath__24_0_in1[9]));
INVX2 inst_cellmath__24_0_I2147 (.Y(N3877), .A(inst_cellmath__24_0_in1[10]));
INVX2 inst_cellmath__24_0_I2155 (.Y(N3885), .A(inst_cellmath__24_0_in1[11]));
INVX1 inst_cellmath__24_0_I2163 (.Y(N3893), .A(inst_cellmath__24_0_in1[12]));
INVX2 inst_cellmath__24_0_I2161 (.Y(N3891), .A(inst_cellmath__24_0_in1[12]));
INVXL inst_cellmath__24_0_I2171 (.Y(N3901), .A(inst_cellmath__24_0_in1[13]));
INVX2 inst_cellmath__24_0_I2170 (.Y(N3900), .A(inst_cellmath__24_0_in1[13]));
INVX3 inst_cellmath__24_0_I2179 (.Y(N3909), .A(inst_cellmath__24_0_in1[14]));
INVX3 inst_cellmath__24_0_I2187 (.Y(N3917), .A(inst_cellmath__24_0_in1[15]));
INVX3 inst_cellmath__24_0_I2195 (.Y(N3925), .A(inst_cellmath__24_0_in1[16]));
INVX3 inst_cellmath__24_0_I2203 (.Y(N3933), .A(inst_cellmath__24_0_in1[17]));
INVX3 inst_cellmath__24_0_I2211 (.Y(N3941), .A(inst_cellmath__24_0_in1[18]));
INVX2 inst_cellmath__24_0_I2219 (.Y(N3949), .A(inst_cellmath__24_0_in1[19]));
INVX3 inst_cellmath__24_0_I2227 (.Y(N3957), .A(inst_cellmath__24_0_in1[20]));
INVX2 inst_cellmath__24_0_I2235 (.Y(N3965), .A(inst_cellmath__24_0_in1[21]));
INVX3 inst_cellmath__24_0_I2243 (.Y(N3973), .A(inst_cellmath__24_0_in1[22]));
INVX1 inst_cellmath__24_0_I2251 (.Y(N3981), .A(inst_cellmath__24_0_in0[0]));
INVX1 inst_cellmath__24_0_I2247 (.Y(N3977), .A(inst_cellmath__24_0_in0[0]));
NOR2XL inst_cellmath__24_0_I87 (.Y(inst_cellmath__24_0_out0[0]), .A(N3981), .B(N3797));
NOR2XL inst_cellmath__24_0_I88 (.Y(N383), .A(N3981), .B(N3805));
NOR2XL inst_cellmath__24_0_I89 (.Y(N385), .A(N3981), .B(N3813));
NOR2XL inst_cellmath__24_0_I90 (.Y(N387), .A(N3981), .B(N3821));
NOR2XL inst_cellmath__24_0_I91 (.Y(N389), .A(N3981), .B(N3829));
NOR2XL inst_cellmath__24_0_I92 (.Y(N391), .A(N3981), .B(N3837));
NOR2XL inst_cellmath__24_0_I93 (.Y(N393), .A(N3981), .B(N3845));
NOR2XL inst_cellmath__24_0_I94 (.Y(N395), .A(N3981), .B(N3853));
NOR2XL inst_cellmath__24_0_I95 (.Y(N397), .A(N3981), .B(N3861));
NOR2XL inst_cellmath__24_0_I96 (.Y(N399), .A(N3981), .B(N3869));
NOR2XL inst_cellmath__24_0_I97 (.Y(N401), .A(N3981), .B(N3877));
NOR2XL inst_cellmath__24_0_I98 (.Y(N403), .A(N3981), .B(N3885));
NOR2XL inst_cellmath__24_0_I99 (.Y(N405), .A(N3981), .B(N3893));
NOR2XL inst_cellmath__24_0_I100 (.Y(N407), .A(N3981), .B(N3901));
NOR2XL inst_cellmath__24_0_I101 (.Y(N409), .A(N3981), .B(N3909));
NOR2XL inst_cellmath__24_0_I102 (.Y(N411), .A(N3981), .B(N3917));
NOR2XL inst_cellmath__24_0_I103 (.Y(N413), .A(N3981), .B(N3925));
NOR2XL inst_cellmath__24_0_I104 (.Y(N415), .A(N3981), .B(N3933));
NOR2XL inst_cellmath__24_0_I105 (.Y(N417), .A(N3981), .B(N3941));
NOR2XL inst_cellmath__24_0_I106 (.Y(N419), .A(N3977), .B(N3949));
NOR2XL inst_cellmath__24_0_I107 (.Y(N421), .A(N3977), .B(N3957));
NOR2XL inst_cellmath__24_0_I108 (.Y(N423), .A(N3977), .B(N3965));
NOR2XL inst_cellmath__24_0_I109 (.Y(N425), .A(N3977), .B(N3973));
INVXL inst_cellmath__24_0_I110 (.Y(N427), .A(N3977));
INVX2 inst_cellmath__24_0_I2259 (.Y(N3989), .A(inst_cellmath__24_0_in0[1]));
NOR2XL inst_cellmath__24_0_I116 (.Y(N440), .A(N3989), .B(N3797));
NOR2XL inst_cellmath__24_0_I117 (.Y(N442), .A(N3989), .B(N3805));
NOR2XL inst_cellmath__24_0_I118 (.Y(N444), .A(N3989), .B(N3813));
NOR2XL inst_cellmath__24_0_I119 (.Y(N446), .A(N3989), .B(N3821));
NOR2XL inst_cellmath__24_0_I120 (.Y(N448), .A(N3989), .B(N3829));
NOR2XL inst_cellmath__24_0_I121 (.Y(N450), .A(N3989), .B(N3837));
NOR2XL inst_cellmath__24_0_I122 (.Y(N452), .A(N3989), .B(N3845));
NOR2XL inst_cellmath__24_0_I123 (.Y(N454), .A(N3989), .B(N3853));
NOR2XL inst_cellmath__24_0_I124 (.Y(N456), .A(N3989), .B(N3861));
NOR2XL inst_cellmath__24_0_I125 (.Y(N458), .A(N3989), .B(N3869));
NOR2XL inst_cellmath__24_0_I126 (.Y(N460), .A(N3989), .B(N3877));
NOR2XL inst_cellmath__24_0_I127 (.Y(N462), .A(N3989), .B(N3885));
NOR2XL inst_cellmath__24_0_I128 (.Y(N464), .A(N3989), .B(N3893));
NOR2XL inst_cellmath__24_0_I129 (.Y(N466), .A(N3989), .B(N3901));
NOR2XL inst_cellmath__24_0_I130 (.Y(N468), .A(N3989), .B(N3909));
NOR2XL inst_cellmath__24_0_I131 (.Y(N470), .A(N3989), .B(N3917));
NOR2XL inst_cellmath__24_0_I132 (.Y(N472), .A(N3989), .B(N3925));
NOR2XL inst_cellmath__24_0_I133 (.Y(N474), .A(N3989), .B(N3933));
NOR2XL inst_cellmath__24_0_I134 (.Y(N476), .A(N3989), .B(N3941));
NOR2X1 inst_cellmath__24_0_I135 (.Y(N478), .A(N3989), .B(N3949));
NOR2XL inst_cellmath__24_0_I136 (.Y(N480), .A(N3989), .B(N3957));
NOR2XL inst_cellmath__24_0_I137 (.Y(N482), .A(N3989), .B(N3965));
NOR2X1 inst_cellmath__24_0_I138 (.Y(N484), .A(N3989), .B(N3973));
INVXL inst_cellmath__24_0_I139 (.Y(N486), .A(N3989));
INVX2 inst_cellmath__24_0_I2267 (.Y(N3997), .A(inst_cellmath__24_0_in0[2]));
INVX3 inst_cellmath__24_0_I2264 (.Y(N3994), .A(inst_cellmath__24_0_in0[2]));
NOR2XL inst_cellmath__24_0_I145 (.Y(N499), .A(N3997), .B(N3797));
NOR2XL inst_cellmath__24_0_I146 (.Y(N501), .A(N3997), .B(N3805));
NOR2XL inst_cellmath__24_0_I147 (.Y(N503), .A(N3997), .B(N3813));
NOR2XL inst_cellmath__24_0_I148 (.Y(N505), .A(N3997), .B(N3821));
NOR2XL inst_cellmath__24_0_I149 (.Y(N507), .A(N3997), .B(N3829));
NOR2XL inst_cellmath__24_0_I150 (.Y(N509), .A(N3997), .B(N3837));
NOR2XL inst_cellmath__24_0_I151 (.Y(N511), .A(N3997), .B(N3845));
NOR2XL inst_cellmath__24_0_I152 (.Y(N513), .A(N3997), .B(N3853));
NOR2XL inst_cellmath__24_0_I153 (.Y(N515), .A(N3997), .B(N3861));
NOR2XL inst_cellmath__24_0_I154 (.Y(N517), .A(N3997), .B(N3869));
NOR2XL inst_cellmath__24_0_I155 (.Y(N519), .A(N3997), .B(N3877));
NOR2X1 inst_cellmath__24_0_I156 (.Y(N521), .A(N3997), .B(N3885));
NOR2XL inst_cellmath__24_0_I157 (.Y(N523), .A(N3997), .B(N3893));
NOR2XL inst_cellmath__24_0_I158 (.Y(N525), .A(N3997), .B(N3901));
NOR2XL inst_cellmath__24_0_I159 (.Y(N527), .A(N3994), .B(N3909));
NOR2X1 inst_cellmath__24_0_I160 (.Y(N529), .A(N3994), .B(N3917));
NOR2XL inst_cellmath__24_0_I161 (.Y(N531), .A(N3994), .B(N3925));
NOR2X1 inst_cellmath__24_0_I162 (.Y(N533), .A(N3994), .B(N3933));
NOR2X1 inst_cellmath__24_0_I163 (.Y(N535), .A(N3994), .B(N3941));
NOR2X1 inst_cellmath__24_0_I164 (.Y(N537), .A(N3994), .B(N3949));
NOR2X1 inst_cellmath__24_0_I165 (.Y(N539), .A(N3994), .B(N3957));
NOR2X2 inst_cellmath__24_0_I166 (.Y(N541), .A(N3994), .B(N3965));
NOR2XL inst_cellmath__24_0_I167 (.Y(N543), .A(N3994), .B(N3973));
INVXL inst_cellmath__24_0_I168 (.Y(N545), .A(N3994));
INVXL inst_cellmath__24_0_I2274 (.Y(N4004), .A(inst_cellmath__24_0_in0[3]));
INVX3 inst_cellmath__24_0_I2273 (.Y(N4003), .A(inst_cellmath__24_0_in0[3]));
NOR2XL inst_cellmath__24_0_I174 (.Y(N558), .A(N4004), .B(N3797));
NOR2XL inst_cellmath__24_0_I175 (.Y(N560), .A(N4004), .B(N3805));
NOR2XL inst_cellmath__24_0_I176 (.Y(N562), .A(N4004), .B(N3813));
NOR2XL inst_cellmath__24_0_I177 (.Y(N564), .A(N4003), .B(N3821));
NOR2XL inst_cellmath__24_0_I178 (.Y(N566), .A(N4003), .B(N3829));
NOR2X2 inst_cellmath__24_0_I179 (.Y(N568), .A(N4003), .B(N3837));
NOR2XL inst_cellmath__24_0_I180 (.Y(N570), .A(N4003), .B(N3845));
NOR2XL inst_cellmath__24_0_I181 (.Y(N572), .A(N4003), .B(N3853));
NOR2XL inst_cellmath__24_0_I182 (.Y(N574), .A(N4003), .B(N3861));
NOR2XL inst_cellmath__24_0_I183 (.Y(N576), .A(N4003), .B(N3869));
NOR2X1 inst_cellmath__24_0_I184 (.Y(N578), .A(N4003), .B(N3877));
NOR2XL inst_cellmath__24_0_I185 (.Y(N580), .A(N4003), .B(N3885));
NOR2XL inst_cellmath__24_0_I186 (.Y(N582), .A(N4003), .B(N3893));
NOR2XL inst_cellmath__24_0_I187 (.Y(N584), .A(N4003), .B(N3901));
NOR2XL inst_cellmath__24_0_I188 (.Y(N586), .A(N4003), .B(N3909));
NOR2XL inst_cellmath__24_0_I189 (.Y(N588), .A(N4003), .B(N3917));
NOR2X1 inst_cellmath__24_0_I190 (.Y(N590), .A(N4003), .B(N3925));
NOR2X2 inst_cellmath__24_0_I191 (.Y(N592), .A(N4003), .B(N3933));
NOR2X1 inst_cellmath__24_0_I192 (.Y(N594), .A(N4003), .B(N3941));
NOR2XL inst_cellmath__24_0_I193 (.Y(N596), .A(N4003), .B(N3949));
NOR2XL inst_cellmath__24_0_I194 (.Y(N598), .A(N4003), .B(N3957));
NOR2X1 inst_cellmath__24_0_I195 (.Y(N600), .A(N4003), .B(N3965));
NOR2XL inst_cellmath__24_0_I196 (.Y(N602), .A(N4003), .B(N3973));
INVXL inst_cellmath__24_0_I197 (.Y(N604), .A(N4003));
INVXL inst_cellmath__24_0_I2281 (.Y(N4011), .A(inst_cellmath__24_0_in0[4]));
INVX2 inst_cellmath__24_0_I2280 (.Y(N4010), .A(inst_cellmath__24_0_in0[4]));
INVX2 inst_cellmath__24_0_I2277 (.Y(N4007), .A(inst_cellmath__24_0_in0[4]));
NOR2XL inst_cellmath__24_0_I203 (.Y(N617), .A(N4011), .B(N3797));
NOR2XL inst_cellmath__24_0_I204 (.Y(N619), .A(N4011), .B(N3805));
NOR2XL inst_cellmath__24_0_I205 (.Y(N621), .A(N4011), .B(N3813));
NOR2XL inst_cellmath__24_0_I206 (.Y(N623), .A(N4011), .B(N3820));
NOR2X2 inst_cellmath__24_0_I207 (.Y(N625), .A(N4010), .B(N3829));
NOR2XL inst_cellmath__24_0_I208 (.Y(N627), .A(N4010), .B(N3837));
NOR2XL inst_cellmath__24_0_I209 (.Y(N629), .A(N4010), .B(N3845));
NOR2XL inst_cellmath__24_0_I210 (.Y(N631), .A(N4010), .B(N3853));
NOR2XL inst_cellmath__24_0_I211 (.Y(N633), .A(N4010), .B(N3861));
NOR2XL inst_cellmath__24_0_I212 (.Y(N635), .A(N4010), .B(N3869));
NOR2XL inst_cellmath__24_0_I213 (.Y(N637), .A(N4010), .B(N3877));
NOR2XL inst_cellmath__24_0_I214 (.Y(N639), .A(N4010), .B(N3885));
NOR2XL inst_cellmath__24_0_I215 (.Y(N641), .A(N4010), .B(N3893));
NOR2X2 inst_cellmath__24_0_I216 (.Y(N643), .A(N4010), .B(N3900));
NOR2XL inst_cellmath__24_0_I217 (.Y(N645), .A(N4010), .B(N3909));
NOR2XL inst_cellmath__24_0_I218 (.Y(N647), .A(N4010), .B(N3917));
NOR2XL inst_cellmath__24_0_I219 (.Y(N649), .A(N4010), .B(N3925));
NOR2XL inst_cellmath__24_0_I220 (.Y(N651), .A(N4010), .B(N3933));
NOR2X1 inst_cellmath__24_0_I221 (.Y(N653), .A(N4010), .B(N3941));
NOR2X1 inst_cellmath__24_0_I222 (.Y(N655), .A(N4007), .B(N3949));
NOR2X1 inst_cellmath__24_0_I223 (.Y(N657), .A(N4007), .B(N3957));
NOR2X2 inst_cellmath__24_0_I224 (.Y(N659), .A(N4007), .B(N3965));
NOR2XL inst_cellmath__24_0_I225 (.Y(N661), .A(N4007), .B(N3973));
INVXL inst_cellmath__24_0_I226 (.Y(N663), .A(N4007));
INVXL inst_cellmath__24_0_I2288 (.Y(N4018), .A(inst_cellmath__24_0_in0[5]));
INVX1 inst_cellmath__24_0_I2287 (.Y(N4017), .A(inst_cellmath__24_0_in0[5]));
INVX3 inst_cellmath__24_0_I2286 (.Y(N4016), .A(inst_cellmath__24_0_in0[5]));
NOR2XL inst_cellmath__24_0_I232 (.Y(N676), .A(N4018), .B(N3797));
NOR2XL inst_cellmath__24_0_I233 (.Y(N678), .A(N4018), .B(N3805));
NOR2XL inst_cellmath__24_0_I234 (.Y(N680), .A(N4018), .B(N3813));
NOR2X1 inst_cellmath__24_0_I235 (.Y(N682), .A(N4017), .B(N3820));
NOR2XL inst_cellmath__24_0_I236 (.Y(N684), .A(N4017), .B(N3829));
NOR2XL inst_cellmath__24_0_I237 (.Y(N686), .A(N4017), .B(N3837));
NOR2XL inst_cellmath__24_0_I238 (.Y(N688), .A(N4017), .B(N3845));
NOR2XL inst_cellmath__24_0_I239 (.Y(N690), .A(N4017), .B(N3853));
NOR2XL inst_cellmath__24_0_I240 (.Y(N692), .A(N4017), .B(N3861));
NOR2XL inst_cellmath__24_0_I241 (.Y(N694), .A(N4017), .B(N3869));
NOR2XL inst_cellmath__24_0_I242 (.Y(N696), .A(N4016), .B(N3877));
NOR2XL inst_cellmath__24_0_I243 (.Y(N698), .A(N4016), .B(N3885));
NOR2X1 inst_cellmath__24_0_I244 (.Y(N700), .A(N4016), .B(N3893));
NOR2XL inst_cellmath__24_0_I245 (.Y(N702), .A(N4016), .B(N3900));
NOR2X1 inst_cellmath__24_0_I246 (.Y(N704), .A(N4016), .B(N3909));
NOR2X2 inst_cellmath__24_0_I247 (.Y(N706), .A(N4016), .B(N3917));
NOR2X1 inst_cellmath__24_0_I248 (.Y(N708), .A(N4016), .B(N3925));
NOR2X1 inst_cellmath__24_0_I249 (.Y(N710), .A(N4016), .B(N3933));
NOR2X1 inst_cellmath__24_0_I250 (.Y(N712), .A(N4016), .B(N3941));
NOR2X2 inst_cellmath__24_0_I251 (.Y(N714), .A(N4016), .B(N3949));
NOR2X1 inst_cellmath__24_0_I252 (.Y(N716), .A(N4016), .B(N3957));
NOR2X1 inst_cellmath__24_0_I253 (.Y(N718), .A(N4016), .B(N3965));
NOR2XL inst_cellmath__24_0_I254 (.Y(N720), .A(N4016), .B(N3973));
INVXL inst_cellmath__24_0_I255 (.Y(N722), .A(N4016));
INVX2 inst_cellmath__24_0_I2295 (.Y(N4025), .A(inst_cellmath__24_0_in0[6]));
INVX2 inst_cellmath__24_0_I2293 (.Y(N4023), .A(inst_cellmath__24_0_in0[6]));
NOR2XL inst_cellmath__24_0_I261 (.Y(N735), .A(N4025), .B(N3797));
NOR2XL inst_cellmath__24_0_I262 (.Y(N737), .A(N4025), .B(N3805));
NOR2X1 inst_cellmath__24_0_I263 (.Y(N739), .A(N4025), .B(N3813));
NOR2XL inst_cellmath__24_0_I264 (.Y(N741), .A(N4025), .B(N3820));
NOR2XL inst_cellmath__24_0_I265 (.Y(N743), .A(N4025), .B(N3829));
NOR2XL inst_cellmath__24_0_I266 (.Y(N745), .A(N4025), .B(N3837));
NOR2XL inst_cellmath__24_0_I267 (.Y(N747), .A(N4025), .B(N3845));
NOR2XL inst_cellmath__24_0_I268 (.Y(N749), .A(N4025), .B(N3853));
NOR2XL inst_cellmath__24_0_I269 (.Y(N751), .A(N4025), .B(N3861));
NOR2XL inst_cellmath__24_0_I270 (.Y(N753), .A(N4023), .B(N3869));
NOR2XL inst_cellmath__24_0_I271 (.Y(N755), .A(N4023), .B(N3877));
NOR2X1 inst_cellmath__24_0_I272 (.Y(N757), .A(N4023), .B(N3885));
NOR2X1 inst_cellmath__24_0_I273 (.Y(N759), .A(N4023), .B(N3893));
NOR2X2 inst_cellmath__24_0_I274 (.Y(N761), .A(N4023), .B(N3900));
NOR2X2 inst_cellmath__24_0_I275 (.Y(N763), .A(N4023), .B(N3909));
NOR2XL inst_cellmath__24_0_I276 (.Y(N765), .A(N4023), .B(N3917));
NOR2XL inst_cellmath__24_0_I277 (.Y(N767), .A(N4023), .B(N3925));
NOR2XL inst_cellmath__24_0_I278 (.Y(N769), .A(N4023), .B(N3933));
NOR2X1 inst_cellmath__24_0_I279 (.Y(N771), .A(N4023), .B(N3941));
NOR2XL inst_cellmath__24_0_I280 (.Y(N773), .A(N4025), .B(N3949));
NOR2X1 inst_cellmath__24_0_I281 (.Y(N775), .A(N4025), .B(N3957));
NOR2X1 inst_cellmath__24_0_I282 (.Y(N777), .A(N4025), .B(N3965));
NOR2XL inst_cellmath__24_0_I283 (.Y(N779), .A(N4025), .B(N3973));
INVXL inst_cellmath__24_0_I284 (.Y(N781), .A(N4025));
INVX1 inst_cellmath__24_0_I2303 (.Y(N4033), .A(inst_cellmath__24_0_in0[7]));
INVX3 inst_cellmath__24_0_I2301 (.Y(N4031), .A(inst_cellmath__24_0_in0[7]));
NOR2XL inst_cellmath__24_0_I290 (.Y(N794), .A(N4033), .B(N3797));
NOR2XL inst_cellmath__24_0_I291 (.Y(N796), .A(N4033), .B(N3805));
NOR2XL inst_cellmath__24_0_I292 (.Y(N798), .A(N4033), .B(N3813));
NOR2XL inst_cellmath__24_0_I293 (.Y(N800), .A(N4033), .B(N3820));
NOR2XL inst_cellmath__24_0_I294 (.Y(N802), .A(N4033), .B(N3829));
NOR2XL inst_cellmath__24_0_I295 (.Y(N804), .A(N4033), .B(N3837));
NOR2XL inst_cellmath__24_0_I296 (.Y(N806), .A(N4033), .B(N3845));
NOR2XL inst_cellmath__24_0_I297 (.Y(N808), .A(N4033), .B(N3853));
NOR2XL inst_cellmath__24_0_I298 (.Y(N810), .A(N4033), .B(N3861));
NOR2XL inst_cellmath__24_0_I299 (.Y(N812), .A(N4031), .B(N3869));
NOR2XL inst_cellmath__24_0_I300 (.Y(N814), .A(N4031), .B(N3877));
NOR2XL inst_cellmath__24_0_I301 (.Y(N816), .A(N4031), .B(N3885));
NOR2X1 inst_cellmath__24_0_I302 (.Y(N818), .A(N4031), .B(N3893));
NOR2X1 inst_cellmath__24_0_I303 (.Y(N820), .A(N4031), .B(N3900));
NOR2X1 inst_cellmath__24_0_I304 (.Y(N822), .A(N4031), .B(N3909));
NOR2X1 inst_cellmath__24_0_I305 (.Y(N824), .A(N4031), .B(N3917));
NOR2X1 inst_cellmath__24_0_I306 (.Y(N826), .A(N4031), .B(N3925));
NOR2XL inst_cellmath__24_0_I307 (.Y(N828), .A(N4031), .B(N3933));
NOR2XL inst_cellmath__24_0_I308 (.Y(N830), .A(N4031), .B(N3941));
NOR2XL inst_cellmath__24_0_I309 (.Y(N832), .A(N4031), .B(N3949));
NOR2XL inst_cellmath__24_0_I310 (.Y(N834), .A(N4031), .B(N3957));
NOR2X1 inst_cellmath__24_0_I311 (.Y(N836), .A(N4031), .B(N3965));
NOR2XL inst_cellmath__24_0_I312 (.Y(N838), .A(N4031), .B(N3973));
INVXL inst_cellmath__24_0_I313 (.Y(N840), .A(N4031));
INVX1 inst_cellmath__24_0_I2311 (.Y(N4041), .A(inst_cellmath__24_0_in0[8]));
INVX3 inst_cellmath__24_0_I2309 (.Y(N4039), .A(inst_cellmath__24_0_in0[8]));
NOR2XL inst_cellmath__24_0_I319 (.Y(N853), .A(N4041), .B(N3797));
NOR2XL inst_cellmath__24_0_I320 (.Y(N855), .A(N4041), .B(N3805));
NOR2XL inst_cellmath__24_0_I321 (.Y(N857), .A(N4041), .B(N3813));
NOR2XL inst_cellmath__24_0_I322 (.Y(N859), .A(N4041), .B(N3820));
NOR2XL inst_cellmath__24_0_I323 (.Y(N861), .A(N4041), .B(N3829));
NOR2XL inst_cellmath__24_0_I324 (.Y(N863), .A(N4041), .B(N3837));
NOR2XL inst_cellmath__24_0_I325 (.Y(N865), .A(N4041), .B(N3845));
NOR2XL inst_cellmath__24_0_I326 (.Y(N867), .A(N4041), .B(N3853));
NOR2XL inst_cellmath__24_0_I327 (.Y(N869), .A(N4041), .B(N3861));
NOR2XL inst_cellmath__24_0_I328 (.Y(N871), .A(N4039), .B(N3869));
NOR2XL inst_cellmath__24_0_I329 (.Y(N873), .A(N4039), .B(N3877));
NOR2X1 inst_cellmath__24_0_I330 (.Y(N875), .A(N4039), .B(N3885));
NOR2X1 inst_cellmath__24_0_I331 (.Y(N877), .A(N4039), .B(N3893));
NOR2X2 inst_cellmath__24_0_I332 (.Y(N879), .A(N4039), .B(N3900));
NOR2XL inst_cellmath__24_0_I333 (.Y(N881), .A(N4039), .B(N3909));
NOR2X1 inst_cellmath__24_0_I334 (.Y(N883), .A(N4039), .B(N3917));
NOR2X1 inst_cellmath__24_0_I335 (.Y(N885), .A(N4039), .B(N3925));
NOR2X1 inst_cellmath__24_0_I336 (.Y(N887), .A(N4039), .B(N3933));
NOR2X1 inst_cellmath__24_0_I337 (.Y(N889), .A(N4039), .B(N3941));
NOR2XL inst_cellmath__24_0_I338 (.Y(N891), .A(N4039), .B(N3949));
NOR2XL inst_cellmath__24_0_I339 (.Y(N893), .A(N4039), .B(N3957));
NOR2XL inst_cellmath__24_0_I340 (.Y(N895), .A(N4039), .B(N3965));
NOR2XL inst_cellmath__24_0_I341 (.Y(N897), .A(N4039), .B(N3973));
INVXL inst_cellmath__24_0_I342 (.Y(N899), .A(N4039));
INVXL inst_cellmath__24_0_I2318 (.Y(N4048), .A(inst_cellmath__24_0_in0[9]));
CLKINVX4 inst_cellmath__24_0_I2317 (.Y(N4047), .A(inst_cellmath__24_0_in0[9]));
NOR2XL inst_cellmath__24_0_I348 (.Y(N912), .A(N4048), .B(N3797));
NOR2XL inst_cellmath__24_0_I349 (.Y(N914), .A(N4048), .B(N3805));
NOR2XL inst_cellmath__24_0_I350 (.Y(N916), .A(N4048), .B(N3813));
NOR2XL inst_cellmath__24_0_I351 (.Y(N918), .A(N4047), .B(N3821));
NOR2XL inst_cellmath__24_0_I352 (.Y(N920), .A(N4047), .B(N3829));
NOR2XL inst_cellmath__24_0_I353 (.Y(N922), .A(N4047), .B(N3837));
NOR2XL inst_cellmath__24_0_I354 (.Y(N924), .A(N4047), .B(N3845));
NOR2XL inst_cellmath__24_0_I355 (.Y(N926), .A(N4047), .B(N3853));
NOR2XL inst_cellmath__24_0_I356 (.Y(N928), .A(N4047), .B(N3861));
NOR2XL inst_cellmath__24_0_I357 (.Y(N930), .A(N4047), .B(N3869));
NOR2XL inst_cellmath__24_0_I358 (.Y(N932), .A(N4047), .B(N3877));
NOR2X2 inst_cellmath__24_0_I359 (.Y(N934), .A(N4047), .B(N3885));
NOR2X1 inst_cellmath__24_0_I360 (.Y(N936), .A(N4047), .B(N3891));
NOR2X2 inst_cellmath__24_0_I361 (.Y(N938), .A(N4047), .B(N3900));
NOR2XL inst_cellmath__24_0_I362 (.Y(N940), .A(N4047), .B(N3909));
NOR2X2 inst_cellmath__24_0_I363 (.Y(N942), .A(N4047), .B(N3917));
NOR2XL inst_cellmath__24_0_I364 (.Y(N944), .A(N4047), .B(N3925));
NOR2X1 inst_cellmath__24_0_I365 (.Y(N946), .A(N4047), .B(N3933));
NOR2XL inst_cellmath__24_0_I366 (.Y(N948), .A(N4047), .B(N3941));
NOR2XL inst_cellmath__24_0_I367 (.Y(N950), .A(N4047), .B(N3949));
NOR2XL inst_cellmath__24_0_I368 (.Y(N952), .A(N4047), .B(N3957));
NOR2XL inst_cellmath__24_0_I369 (.Y(N954), .A(N4047), .B(N3965));
NOR2XL inst_cellmath__24_0_I370 (.Y(N956), .A(N4047), .B(N3973));
INVXL inst_cellmath__24_0_I371 (.Y(N958), .A(N4047));
INVXL inst_cellmath__24_0_I2325 (.Y(N4055), .A(inst_cellmath__24_0_in0[10]));
INVX3 inst_cellmath__24_0_I2323 (.Y(N4053), .A(inst_cellmath__24_0_in0[10]));
NOR2XL inst_cellmath__24_0_I377 (.Y(N971), .A(N4055), .B(N3797));
NOR2XL inst_cellmath__24_0_I378 (.Y(N973), .A(N4055), .B(N3805));
NOR2XL inst_cellmath__24_0_I379 (.Y(N975), .A(N4055), .B(N3813));
NOR2XL inst_cellmath__24_0_I380 (.Y(N977), .A(N4055), .B(N3821));
NOR2XL inst_cellmath__24_0_I381 (.Y(N979), .A(N4055), .B(N3829));
NOR2XL inst_cellmath__24_0_I382 (.Y(N981), .A(N4055), .B(N3837));
NOR2XL inst_cellmath__24_0_I383 (.Y(N983), .A(N4055), .B(N3845));
NOR2XL inst_cellmath__24_0_I384 (.Y(N985), .A(N4055), .B(N3853));
NOR2XL inst_cellmath__24_0_I385 (.Y(N987), .A(N4055), .B(N3861));
NOR2XL inst_cellmath__24_0_I386 (.Y(N989), .A(N4053), .B(N3869));
NOR2XL inst_cellmath__24_0_I387 (.Y(N991), .A(N4053), .B(N3877));
NOR2X1 inst_cellmath__24_0_I388 (.Y(N993), .A(N4053), .B(N3885));
NOR2X1 inst_cellmath__24_0_I389 (.Y(N995), .A(N4053), .B(N3891));
NOR2X1 inst_cellmath__24_0_I390 (.Y(N997), .A(N4053), .B(N3900));
NOR2XL inst_cellmath__24_0_I391 (.Y(N999), .A(N4053), .B(N3909));
NOR2X1 inst_cellmath__24_0_I392 (.Y(N1001), .A(N4053), .B(N3917));
NOR2XL inst_cellmath__24_0_I393 (.Y(N1003), .A(N4053), .B(N3925));
NOR2XL inst_cellmath__24_0_I394 (.Y(N1005), .A(N4053), .B(N3933));
NOR2XL inst_cellmath__24_0_I395 (.Y(N1007), .A(N4053), .B(N3941));
NOR2XL inst_cellmath__24_0_I396 (.Y(N1009), .A(N4053), .B(N3949));
NOR2XL inst_cellmath__24_0_I397 (.Y(N1011), .A(N4053), .B(N3957));
NOR2XL inst_cellmath__24_0_I398 (.Y(N1013), .A(N4053), .B(N3965));
NOR2XL inst_cellmath__24_0_I399 (.Y(N1015), .A(N4053), .B(N3973));
INVXL inst_cellmath__24_0_I400 (.Y(N1017), .A(N4053));
CLKINVX4 inst_cellmath__24_0_I2333 (.Y(N4063), .A(inst_cellmath__24_0_in0[11]));
NOR2XL inst_cellmath__24_0_I406 (.Y(N1030), .A(N4063), .B(N3797));
NOR2XL inst_cellmath__24_0_I407 (.Y(N1032), .A(N4063), .B(N3805));
NOR2XL inst_cellmath__24_0_I408 (.Y(N1034), .A(N4063), .B(N3813));
NOR2XL inst_cellmath__24_0_I409 (.Y(N1036), .A(N4063), .B(N3821));
NOR2XL inst_cellmath__24_0_I410 (.Y(N1038), .A(N4063), .B(N3829));
NOR2XL inst_cellmath__24_0_I411 (.Y(N1040), .A(N4063), .B(N3837));
NOR2XL inst_cellmath__24_0_I412 (.Y(N1042), .A(N4063), .B(N3845));
NOR2XL inst_cellmath__24_0_I413 (.Y(N1044), .A(N4063), .B(N3853));
NOR2X1 inst_cellmath__24_0_I414 (.Y(N1046), .A(N4063), .B(N3861));
NOR2XL inst_cellmath__24_0_I415 (.Y(N1048), .A(N4063), .B(N3869));
NOR2X1 inst_cellmath__24_0_I416 (.Y(N1050), .A(N4063), .B(N3877));
NOR2XL inst_cellmath__24_0_I417 (.Y(N1052), .A(N4063), .B(N3885));
NOR2X1 inst_cellmath__24_0_I418 (.Y(N1054), .A(N4063), .B(N3891));
NOR2X1 inst_cellmath__24_0_I419 (.Y(N1056), .A(N4063), .B(N3900));
NOR2X1 inst_cellmath__24_0_I420 (.Y(N1058), .A(N4063), .B(N3909));
NOR2XL inst_cellmath__24_0_I421 (.Y(N1060), .A(N4063), .B(N3917));
NOR2XL inst_cellmath__24_0_I422 (.Y(N1062), .A(N4063), .B(N3925));
NOR2XL inst_cellmath__24_0_I423 (.Y(N1064), .A(N4063), .B(N3933));
NOR2XL inst_cellmath__24_0_I424 (.Y(N1066), .A(N4063), .B(N3941));
NOR2XL inst_cellmath__24_0_I425 (.Y(N1068), .A(N4063), .B(N3949));
NOR2XL inst_cellmath__24_0_I426 (.Y(N1070), .A(N4063), .B(N3957));
NOR2XL inst_cellmath__24_0_I427 (.Y(N1072), .A(N4063), .B(N3965));
NOR2XL inst_cellmath__24_0_I428 (.Y(N1074), .A(N4063), .B(N3973));
INVXL inst_cellmath__24_0_I429 (.Y(N1076), .A(N4063));
INVXL inst_cellmath__24_0_I2341 (.Y(N4071), .A(inst_cellmath__24_0_in0[12]));
INVX2 inst_cellmath__24_0_I2340 (.Y(N4070), .A(inst_cellmath__24_0_in0[12]));
INVX2 inst_cellmath__24_0_I2338 (.Y(N4068), .A(inst_cellmath__24_0_in0[12]));
NOR2XL inst_cellmath__24_0_I435 (.Y(N1089), .A(N4071), .B(N3797));
NOR2XL inst_cellmath__24_0_I436 (.Y(N1091), .A(N4071), .B(N3805));
NOR2XL inst_cellmath__24_0_I437 (.Y(N1093), .A(N4071), .B(N3813));
NOR2XL inst_cellmath__24_0_I438 (.Y(N1095), .A(N4071), .B(N3821));
NOR2XL inst_cellmath__24_0_I439 (.Y(N1097), .A(N4070), .B(N3829));
NOR2XL inst_cellmath__24_0_I440 (.Y(N1099), .A(N4070), .B(N3837));
NOR2XL inst_cellmath__24_0_I441 (.Y(N1101), .A(N4070), .B(N3845));
NOR2X1 inst_cellmath__24_0_I442 (.Y(N1103), .A(N4070), .B(N3853));
NOR2XL inst_cellmath__24_0_I443 (.Y(N1105), .A(N4070), .B(N3861));
NOR2X1 inst_cellmath__24_0_I444 (.Y(N1107), .A(N4070), .B(N3869));
NOR2XL inst_cellmath__24_0_I445 (.Y(N1109), .A(N4070), .B(N3877));
NOR2XL inst_cellmath__24_0_I446 (.Y(N1111), .A(N4070), .B(N3885));
NOR2X1 inst_cellmath__24_0_I447 (.Y(N1113), .A(N4070), .B(N3891));
NOR2XL inst_cellmath__24_0_I448 (.Y(N1115), .A(N4070), .B(N3900));
NOR2XL inst_cellmath__24_0_I449 (.Y(N1117), .A(N4068), .B(N3909));
NOR2XL inst_cellmath__24_0_I450 (.Y(N1119), .A(N4068), .B(N3917));
NOR2XL inst_cellmath__24_0_I451 (.Y(N1121), .A(N4068), .B(N3925));
NOR2XL inst_cellmath__24_0_I452 (.Y(N1123), .A(N4068), .B(N3933));
NOR2XL inst_cellmath__24_0_I453 (.Y(N1125), .A(N4068), .B(N3941));
NOR2XL inst_cellmath__24_0_I454 (.Y(N1127), .A(N4068), .B(N3949));
NOR2XL inst_cellmath__24_0_I455 (.Y(N1129), .A(N4068), .B(N3957));
NOR2XL inst_cellmath__24_0_I456 (.Y(N1131), .A(N4068), .B(N3965));
NOR2XL inst_cellmath__24_0_I457 (.Y(N1133), .A(N4068), .B(N3973));
INVXL inst_cellmath__24_0_I458 (.Y(N1135), .A(N4068));
INVXL inst_cellmath__24_0_I2349 (.Y(N4079), .A(inst_cellmath__24_0_in0[13]));
INVX3 inst_cellmath__24_0_I2348 (.Y(N4078), .A(inst_cellmath__24_0_in0[13]));
NOR2XL inst_cellmath__24_0_I464 (.Y(N1148), .A(N4079), .B(N3797));
NOR2XL inst_cellmath__24_0_I465 (.Y(N1150), .A(N4079), .B(N3805));
NOR2XL inst_cellmath__24_0_I466 (.Y(N1152), .A(N4079), .B(N3813));
NOR2XL inst_cellmath__24_0_I467 (.Y(N1154), .A(N4079), .B(N3821));
NOR2XL inst_cellmath__24_0_I468 (.Y(N1156), .A(N4078), .B(N3829));
NOR2XL inst_cellmath__24_0_I469 (.Y(N1158), .A(N4078), .B(N3837));
NOR2XL inst_cellmath__24_0_I470 (.Y(N1160), .A(N4078), .B(N3845));
NOR2XL inst_cellmath__24_0_I471 (.Y(N1162), .A(N4078), .B(N3853));
NOR2XL inst_cellmath__24_0_I472 (.Y(N1164), .A(N4078), .B(N3861));
NOR2XL inst_cellmath__24_0_I473 (.Y(N1166), .A(N4078), .B(N3869));
NOR2X1 inst_cellmath__24_0_I474 (.Y(N1168), .A(N4078), .B(N3877));
NOR2XL inst_cellmath__24_0_I475 (.Y(N1170), .A(N4078), .B(N3885));
NOR2X1 inst_cellmath__24_0_I476 (.Y(N1172), .A(N4078), .B(N3891));
NOR2XL inst_cellmath__24_0_I477 (.Y(N1174), .A(N4078), .B(N3900));
NOR2XL inst_cellmath__24_0_I478 (.Y(N1176), .A(N4078), .B(N3909));
NOR2XL inst_cellmath__24_0_I479 (.Y(N1178), .A(N4078), .B(N3917));
NOR2XL inst_cellmath__24_0_I480 (.Y(N1180), .A(N4078), .B(N3925));
NOR2XL inst_cellmath__24_0_I481 (.Y(N1182), .A(N4078), .B(N3933));
NOR2XL inst_cellmath__24_0_I482 (.Y(N1184), .A(N4078), .B(N3941));
NOR2XL inst_cellmath__24_0_I483 (.Y(N1186), .A(N4078), .B(N3949));
NOR2XL inst_cellmath__24_0_I484 (.Y(N1188), .A(N4078), .B(N3957));
NOR2XL inst_cellmath__24_0_I485 (.Y(N1190), .A(N4078), .B(N3965));
NOR2XL inst_cellmath__24_0_I486 (.Y(N1192), .A(N4078), .B(N3973));
INVXL inst_cellmath__24_0_I487 (.Y(N1194), .A(N4078));
CLKINVX4 inst_cellmath__24_0_I2357 (.Y(N4087), .A(inst_cellmath__24_0_in0[14]));
NOR2XL inst_cellmath__24_0_I493 (.Y(N1207), .A(N4087), .B(N3797));
NOR2XL inst_cellmath__24_0_I494 (.Y(N1209), .A(N4087), .B(N3805));
NOR2XL inst_cellmath__24_0_I495 (.Y(N1211), .A(N4087), .B(N3813));
NOR2XL inst_cellmath__24_0_I496 (.Y(N1213), .A(N4087), .B(N3820));
NOR2XL inst_cellmath__24_0_I497 (.Y(N1215), .A(N4087), .B(N3826));
NOR2X1 inst_cellmath__24_0_I498 (.Y(N1217), .A(N4087), .B(N3834));
NOR2XL inst_cellmath__24_0_I499 (.Y(N1219), .A(N4087), .B(N3845));
NOR2XL inst_cellmath__24_0_I500 (.Y(N1221), .A(N4087), .B(N3853));
NOR2XL inst_cellmath__24_0_I501 (.Y(N1223), .A(N4087), .B(N3861));
NOR2X1 inst_cellmath__24_0_I502 (.Y(N1225), .A(N4087), .B(N3869));
NOR2X1 inst_cellmath__24_0_I503 (.Y(N1227), .A(N4087), .B(N3877));
NOR2X2 inst_cellmath__24_0_I504 (.Y(N1229), .A(N4087), .B(N3885));
NOR2XL inst_cellmath__24_0_I505 (.Y(N1231), .A(N4087), .B(N3891));
NOR2XL inst_cellmath__24_0_I506 (.Y(N1233), .A(N4087), .B(N3900));
NOR2XL inst_cellmath__24_0_I507 (.Y(N1235), .A(N4087), .B(N3909));
NOR2XL inst_cellmath__24_0_I508 (.Y(N1237), .A(N4087), .B(N3917));
NOR2XL inst_cellmath__24_0_I509 (.Y(N1239), .A(N4087), .B(N3925));
NOR2XL inst_cellmath__24_0_I510 (.Y(N1241), .A(N4087), .B(N3933));
NOR2XL inst_cellmath__24_0_I511 (.Y(N1243), .A(N4087), .B(N3941));
NOR2XL inst_cellmath__24_0_I512 (.Y(N1245), .A(N4087), .B(N3949));
NOR2XL inst_cellmath__24_0_I513 (.Y(N1247), .A(N4087), .B(N3957));
NOR2XL inst_cellmath__24_0_I514 (.Y(N1249), .A(N4087), .B(N3965));
NOR2XL inst_cellmath__24_0_I515 (.Y(N1251), .A(N4087), .B(N3973));
INVXL inst_cellmath__24_0_I516 (.Y(N1253), .A(N4087));
INVX3 inst_cellmath__24_0_I2364 (.Y(N4094), .A(inst_cellmath__24_0_in0[15]));
NOR2XL inst_cellmath__24_0_I522 (.Y(N1266), .A(N4094), .B(N3797));
NOR2XL inst_cellmath__24_0_I523 (.Y(N1268), .A(N4094), .B(N3805));
NOR2XL inst_cellmath__24_0_I524 (.Y(N1270), .A(N4094), .B(N3813));
NOR2XL inst_cellmath__24_0_I525 (.Y(N1272), .A(N4094), .B(N3820));
NOR2X1 inst_cellmath__24_0_I526 (.Y(N1274), .A(N4094), .B(N3826));
NOR2XL inst_cellmath__24_0_I527 (.Y(N1276), .A(N4094), .B(N3834));
NOR2X1 inst_cellmath__24_0_I528 (.Y(N1278), .A(N4094), .B(N3845));
NOR2X1 inst_cellmath__24_0_I529 (.Y(N1280), .A(N4094), .B(N3853));
NOR2XL inst_cellmath__24_0_I530 (.Y(N1282), .A(N4094), .B(N3861));
NOR2X1 inst_cellmath__24_0_I531 (.Y(N1284), .A(N4094), .B(N3869));
NOR2XL inst_cellmath__24_0_I532 (.Y(N1286), .A(N4094), .B(N3877));
NOR2X1 inst_cellmath__24_0_I533 (.Y(N1288), .A(N4094), .B(N3885));
NOR2XL inst_cellmath__24_0_I534 (.Y(N1290), .A(N4094), .B(N3891));
NOR2XL inst_cellmath__24_0_I535 (.Y(N1292), .A(N4094), .B(N3900));
NOR2XL inst_cellmath__24_0_I536 (.Y(N1294), .A(N4094), .B(N3909));
NOR2XL inst_cellmath__24_0_I537 (.Y(N1296), .A(N4094), .B(N3917));
NOR2XL inst_cellmath__24_0_I538 (.Y(N1298), .A(N4094), .B(N3925));
NOR2XL inst_cellmath__24_0_I539 (.Y(N1300), .A(N4094), .B(N3933));
NOR2XL inst_cellmath__24_0_I540 (.Y(N1302), .A(N4094), .B(N3941));
NOR2XL inst_cellmath__24_0_I541 (.Y(N1304), .A(N4094), .B(N3949));
NOR2XL inst_cellmath__24_0_I542 (.Y(N1306), .A(N4094), .B(N3957));
NOR2XL inst_cellmath__24_0_I543 (.Y(N1308), .A(N4094), .B(N3965));
NOR2XL inst_cellmath__24_0_I544 (.Y(N1310), .A(N4094), .B(N3973));
INVXL inst_cellmath__24_0_I545 (.Y(N1312), .A(N4094));
INVX3 inst_cellmath__24_0_I2371 (.Y(N4101), .A(inst_cellmath__24_0_in0[16]));
NOR2XL inst_cellmath__24_0_I551 (.Y(N1325), .A(N4101), .B(N3797));
NOR2XL inst_cellmath__24_0_I552 (.Y(N1327), .A(N4101), .B(N3805));
NOR2XL inst_cellmath__24_0_I553 (.Y(N1329), .A(N4101), .B(N3813));
NOR2XL inst_cellmath__24_0_I554 (.Y(N1331), .A(N4101), .B(N3820));
NOR2XL inst_cellmath__24_0_I555 (.Y(N1333), .A(N4101), .B(N3826));
NOR2XL inst_cellmath__24_0_I556 (.Y(N1335), .A(N4101), .B(N3834));
NOR2X1 inst_cellmath__24_0_I557 (.Y(N1337), .A(N4101), .B(N3845));
NOR2X1 inst_cellmath__24_0_I558 (.Y(N1339), .A(N4101), .B(N3853));
NOR2XL inst_cellmath__24_0_I559 (.Y(N1341), .A(N4101), .B(N3861));
NOR2X1 inst_cellmath__24_0_I560 (.Y(N1343), .A(N4101), .B(N3869));
NOR2XL inst_cellmath__24_0_I561 (.Y(N1345), .A(N4101), .B(N3877));
NOR2X1 inst_cellmath__24_0_I562 (.Y(N1347), .A(N4101), .B(N3885));
NOR2XL inst_cellmath__24_0_I563 (.Y(N1349), .A(N4101), .B(N3891));
NOR2XL inst_cellmath__24_0_I564 (.Y(N1351), .A(N4101), .B(N3900));
NOR2XL inst_cellmath__24_0_I565 (.Y(N1353), .A(N4101), .B(N3909));
NOR2XL inst_cellmath__24_0_I566 (.Y(N1355), .A(N4101), .B(N3917));
NOR2XL inst_cellmath__24_0_I567 (.Y(N1357), .A(N4101), .B(N3925));
NOR2XL inst_cellmath__24_0_I568 (.Y(N1359), .A(N4101), .B(N3933));
NOR2XL inst_cellmath__24_0_I569 (.Y(N1361), .A(N4101), .B(N3941));
NOR2XL inst_cellmath__24_0_I570 (.Y(N1363), .A(N4101), .B(N3949));
NOR2XL inst_cellmath__24_0_I571 (.Y(N1365), .A(N4101), .B(N3957));
NOR2XL inst_cellmath__24_0_I572 (.Y(N1367), .A(N4101), .B(N3965));
NOR2XL inst_cellmath__24_0_I573 (.Y(N1369), .A(N4101), .B(N3973));
INVXL inst_cellmath__24_0_I574 (.Y(N1371), .A(N4101));
INVX3 inst_cellmath__24_0_I2379 (.Y(N4109), .A(inst_cellmath__24_0_in0[17]));
NOR2XL inst_cellmath__24_0_I580 (.Y(N1384), .A(N4109), .B(N3797));
NOR2XL inst_cellmath__24_0_I581 (.Y(N1386), .A(N4109), .B(N3805));
NOR2XL inst_cellmath__24_0_I582 (.Y(N1388), .A(N4109), .B(N3813));
NOR2XL inst_cellmath__24_0_I583 (.Y(N1390), .A(N4109), .B(N3820));
NOR2XL inst_cellmath__24_0_I584 (.Y(N1392), .A(N4109), .B(N3826));
NOR2XL inst_cellmath__24_0_I585 (.Y(N1394), .A(N4109), .B(N3834));
NOR2X1 inst_cellmath__24_0_I586 (.Y(N1396), .A(N4109), .B(N3845));
NOR2X1 inst_cellmath__24_0_I587 (.Y(N1398), .A(N4109), .B(N3853));
NOR2X1 inst_cellmath__24_0_I588 (.Y(N1400), .A(N4109), .B(N3861));
NOR2XL inst_cellmath__24_0_I589 (.Y(N1402), .A(N4109), .B(N3869));
NOR2XL inst_cellmath__24_0_I590 (.Y(N1404), .A(N4109), .B(N3877));
NOR2X1 inst_cellmath__24_0_I591 (.Y(N1406), .A(N4109), .B(N3885));
NOR2XL inst_cellmath__24_0_I592 (.Y(N1408), .A(N4109), .B(N3891));
NOR2XL inst_cellmath__24_0_I593 (.Y(N1410), .A(N4109), .B(N3900));
NOR2XL inst_cellmath__24_0_I594 (.Y(N1412), .A(N4109), .B(N3909));
NOR2XL inst_cellmath__24_0_I595 (.Y(N1414), .A(N4109), .B(N3917));
NOR2XL inst_cellmath__24_0_I596 (.Y(N1416), .A(N4109), .B(N3925));
NOR2XL inst_cellmath__24_0_I597 (.Y(N1418), .A(N4109), .B(N3933));
NOR2XL inst_cellmath__24_0_I598 (.Y(N1420), .A(N4109), .B(N3941));
NOR2XL inst_cellmath__24_0_I599 (.Y(N1422), .A(N4109), .B(N3949));
NOR2XL inst_cellmath__24_0_I600 (.Y(N1424), .A(N4109), .B(N3957));
NOR2XL inst_cellmath__24_0_I601 (.Y(N1426), .A(N4109), .B(N3965));
NOR2XL inst_cellmath__24_0_I602 (.Y(N1428), .A(N4109), .B(N3973));
INVXL inst_cellmath__24_0_I603 (.Y(N1430), .A(N4109));
INVX1 inst_cellmath__24_0_I2387 (.Y(N4117), .A(inst_cellmath__24_0_in0[18]));
INVX2 inst_cellmath__24_0_I2386 (.Y(N4116), .A(inst_cellmath__24_0_in0[18]));
NOR2XL inst_cellmath__24_0_I609 (.Y(N1443), .A(N4117), .B(N3797));
NOR2XL inst_cellmath__24_0_I610 (.Y(N1445), .A(N4117), .B(N3805));
NOR2XL inst_cellmath__24_0_I611 (.Y(N1447), .A(N4117), .B(N3813));
NOR2XL inst_cellmath__24_0_I612 (.Y(N1449), .A(N4117), .B(N3820));
NOR2X1 inst_cellmath__24_0_I613 (.Y(N1451), .A(N4116), .B(N3826));
NOR2XL inst_cellmath__24_0_I614 (.Y(N1453), .A(N4116), .B(N3834));
NOR2X1 inst_cellmath__24_0_I615 (.Y(N1455), .A(N4116), .B(N3845));
NOR2XL inst_cellmath__24_0_I616 (.Y(N1457), .A(N4116), .B(N3853));
NOR2XL inst_cellmath__24_0_I617 (.Y(N1459), .A(N4116), .B(N3861));
NOR2XL inst_cellmath__24_0_I618 (.Y(N1461), .A(N4116), .B(N3869));
NOR2XL inst_cellmath__24_0_I619 (.Y(N1463), .A(N4116), .B(N3877));
NOR2XL inst_cellmath__24_0_I620 (.Y(N1465), .A(N4116), .B(N3885));
NOR2XL inst_cellmath__24_0_I621 (.Y(N1467), .A(N4116), .B(N3891));
NOR2XL inst_cellmath__24_0_I622 (.Y(N1469), .A(N4116), .B(N3900));
NOR2XL inst_cellmath__24_0_I623 (.Y(N1471), .A(N4116), .B(N3909));
NOR2XL inst_cellmath__24_0_I624 (.Y(N1473), .A(N4116), .B(N3917));
NOR2XL inst_cellmath__24_0_I625 (.Y(N1475), .A(N4116), .B(N3925));
NOR2XL inst_cellmath__24_0_I626 (.Y(N1477), .A(N4116), .B(N3933));
NOR2XL inst_cellmath__24_0_I627 (.Y(N1479), .A(N4116), .B(N3941));
NOR2XL inst_cellmath__24_0_I628 (.Y(N1481), .A(N4117), .B(N3949));
NOR2XL inst_cellmath__24_0_I629 (.Y(N1483), .A(N4117), .B(N3957));
NOR2XL inst_cellmath__24_0_I630 (.Y(N1485), .A(N4117), .B(N3965));
NOR2XL inst_cellmath__24_0_I631 (.Y(N1487), .A(N4117), .B(N3973));
INVXL inst_cellmath__24_0_I632 (.Y(N1489), .A(N4117));
INVX2 inst_cellmath__24_0_I2395 (.Y(N4125), .A(inst_cellmath__24_0_in0[19]));
NOR2XL inst_cellmath__24_0_I638 (.Y(N1502), .A(N4125), .B(N3793));
NOR2XL inst_cellmath__24_0_I639 (.Y(N1504), .A(N4125), .B(N3805));
NOR2XL inst_cellmath__24_0_I640 (.Y(N1506), .A(N4125), .B(N3813));
NOR2X1 inst_cellmath__24_0_I641 (.Y(N1508), .A(N4125), .B(N3820));
NOR2X1 inst_cellmath__24_0_I642 (.Y(N1510), .A(N4125), .B(N3826));
NOR2X1 inst_cellmath__24_0_I643 (.Y(N1512), .A(N4125), .B(N3834));
NOR2XL inst_cellmath__24_0_I644 (.Y(N1514), .A(N4125), .B(N3845));
NOR2XL inst_cellmath__24_0_I645 (.Y(N1516), .A(N4125), .B(N3853));
NOR2XL inst_cellmath__24_0_I646 (.Y(N1518), .A(N4125), .B(N3861));
NOR2XL inst_cellmath__24_0_I647 (.Y(N1520), .A(N4125), .B(N3869));
NOR2XL inst_cellmath__24_0_I648 (.Y(N1522), .A(N4125), .B(N3877));
NOR2XL inst_cellmath__24_0_I649 (.Y(N1524), .A(N4125), .B(N3885));
NOR2XL inst_cellmath__24_0_I650 (.Y(N1526), .A(N4125), .B(N3893));
NOR2XL inst_cellmath__24_0_I651 (.Y(N1528), .A(N4125), .B(N3901));
NOR2XL inst_cellmath__24_0_I652 (.Y(N1530), .A(N4125), .B(N3909));
NOR2XL inst_cellmath__24_0_I653 (.Y(N1532), .A(N4125), .B(N3917));
NOR2XL inst_cellmath__24_0_I654 (.Y(N1534), .A(N4125), .B(N3925));
NOR2XL inst_cellmath__24_0_I655 (.Y(N1536), .A(N4125), .B(N3933));
NOR2XL inst_cellmath__24_0_I656 (.Y(N1538), .A(N4125), .B(N3941));
NOR2XL inst_cellmath__24_0_I657 (.Y(N1540), .A(N4125), .B(N3949));
NOR2XL inst_cellmath__24_0_I658 (.Y(N1542), .A(N4125), .B(N3957));
NOR2XL inst_cellmath__24_0_I659 (.Y(N1544), .A(N4125), .B(N3965));
NOR2XL inst_cellmath__24_0_I660 (.Y(N1546), .A(N4125), .B(N3973));
INVXL inst_cellmath__24_0_I661 (.Y(N1548), .A(N4125));
INVX2 inst_cellmath__24_0_I2403 (.Y(N4133), .A(inst_cellmath__24_0_in0[20]));
NOR2XL inst_cellmath__24_0_I667 (.Y(N1561), .A(N4133), .B(N3793));
NOR2XL inst_cellmath__24_0_I668 (.Y(N1563), .A(N4133), .B(N3805));
NOR2XL inst_cellmath__24_0_I669 (.Y(N1565), .A(N4133), .B(N3813));
NOR2X1 inst_cellmath__24_0_I670 (.Y(N1567), .A(N4133), .B(N3820));
NOR2X1 inst_cellmath__24_0_I671 (.Y(N1569), .A(N4133), .B(N3826));
NOR2X1 inst_cellmath__24_0_I672 (.Y(N1571), .A(N4133), .B(N3834));
NOR2XL inst_cellmath__24_0_I673 (.Y(N1573), .A(N4133), .B(N3845));
NOR2XL inst_cellmath__24_0_I674 (.Y(N1575), .A(N4133), .B(N3853));
NOR2XL inst_cellmath__24_0_I675 (.Y(N1577), .A(N4133), .B(N3861));
NOR2XL inst_cellmath__24_0_I676 (.Y(N1579), .A(N4133), .B(N3869));
NOR2XL inst_cellmath__24_0_I677 (.Y(N1581), .A(N4133), .B(N3877));
NOR2XL inst_cellmath__24_0_I678 (.Y(N1583), .A(N4133), .B(N3885));
NOR2XL inst_cellmath__24_0_I679 (.Y(N1585), .A(N4133), .B(N3893));
NOR2XL inst_cellmath__24_0_I680 (.Y(N1587), .A(N4133), .B(N3901));
NOR2XL inst_cellmath__24_0_I681 (.Y(N1589), .A(N4133), .B(N3909));
NOR2XL inst_cellmath__24_0_I682 (.Y(N1591), .A(N4133), .B(N3917));
NOR2XL inst_cellmath__24_0_I683 (.Y(N1593), .A(N4133), .B(N3925));
NOR2XL inst_cellmath__24_0_I684 (.Y(N1595), .A(N4133), .B(N3933));
NOR2XL inst_cellmath__24_0_I685 (.Y(N1597), .A(N4133), .B(N3941));
NOR2XL inst_cellmath__24_0_I686 (.Y(N1599), .A(N4133), .B(N3949));
NOR2XL inst_cellmath__24_0_I687 (.Y(N1601), .A(N4133), .B(N3957));
NOR2XL inst_cellmath__24_0_I688 (.Y(N1603), .A(N4133), .B(N3965));
NOR2XL inst_cellmath__24_0_I689 (.Y(N1605), .A(N4133), .B(N3973));
INVXL inst_cellmath__24_0_I690 (.Y(N1607), .A(N4133));
INVX2 inst_cellmath__24_0_I2411 (.Y(N4141), .A(inst_cellmath__24_0_in0[21]));
NOR2XL inst_cellmath__24_0_I696 (.Y(N1620), .A(N4141), .B(N3793));
NOR2XL inst_cellmath__24_0_I697 (.Y(N1622), .A(N4141), .B(N3805));
NOR2XL inst_cellmath__24_0_I698 (.Y(N1624), .A(N4141), .B(N3813));
NOR2X1 inst_cellmath__24_0_I699 (.Y(N1626), .A(N4141), .B(N3820));
NOR2XL inst_cellmath__24_0_I700 (.Y(N1628), .A(N4141), .B(N3826));
NOR2X1 inst_cellmath__24_0_I701 (.Y(N1630), .A(N4141), .B(N3834));
NOR2XL inst_cellmath__24_0_I702 (.Y(N1632), .A(N4141), .B(N3845));
NOR2XL inst_cellmath__24_0_I703 (.Y(N1634), .A(N4141), .B(N3853));
NOR2XL inst_cellmath__24_0_I704 (.Y(N1636), .A(N4141), .B(N3861));
NOR2XL inst_cellmath__24_0_I705 (.Y(N1638), .A(N4141), .B(N3869));
NOR2XL inst_cellmath__24_0_I706 (.Y(N1640), .A(N4141), .B(N3877));
NOR2XL inst_cellmath__24_0_I707 (.Y(N1642), .A(N4141), .B(N3885));
NOR2XL inst_cellmath__24_0_I708 (.Y(N1644), .A(N4141), .B(N3893));
NOR2XL inst_cellmath__24_0_I709 (.Y(N1646), .A(N4141), .B(N3901));
NOR2XL inst_cellmath__24_0_I710 (.Y(N1648), .A(N4141), .B(N3909));
NOR2XL inst_cellmath__24_0_I711 (.Y(N1650), .A(N4141), .B(N3917));
NOR2XL inst_cellmath__24_0_I712 (.Y(N1652), .A(N4141), .B(N3925));
NOR2XL inst_cellmath__24_0_I713 (.Y(N1654), .A(N4141), .B(N3933));
NOR2XL inst_cellmath__24_0_I714 (.Y(N1656), .A(N4141), .B(N3941));
NOR2XL inst_cellmath__24_0_I715 (.Y(N1658), .A(N4141), .B(N3949));
NOR2XL inst_cellmath__24_0_I716 (.Y(N1660), .A(N4141), .B(N3957));
NOR2XL inst_cellmath__24_0_I717 (.Y(N1662), .A(N4141), .B(N3965));
NOR2XL inst_cellmath__24_0_I718 (.Y(N1664), .A(N4141), .B(N3973));
INVXL inst_cellmath__24_0_I719 (.Y(N1666), .A(N4141));
INVX2 inst_cellmath__24_0_I2884 (.Y(N4149), .A(inst_cellmath__24_0_in0[22]));
NOR2XL inst_cellmath__24_0_I725 (.Y(N1679), .A(N4149), .B(N3793));
NOR2XL inst_cellmath__24_0_I726 (.Y(N1681), .A(N4149), .B(N3805));
NOR2XL inst_cellmath__24_0_I727 (.Y(N1683), .A(N4149), .B(N3813));
NOR2XL inst_cellmath__24_0_I728 (.Y(N1685), .A(N4149), .B(N3820));
NOR2XL inst_cellmath__24_0_I729 (.Y(N1687), .A(N4149), .B(N3826));
NOR2XL inst_cellmath__24_0_I730 (.Y(N1689), .A(N4149), .B(N3834));
NOR2XL inst_cellmath__24_0_I731 (.Y(N1691), .A(N4149), .B(N3845));
NOR2XL inst_cellmath__24_0_I732 (.Y(N1693), .A(N4149), .B(N3853));
NOR2XL inst_cellmath__24_0_I733 (.Y(N1695), .A(N4149), .B(N3861));
NOR2XL inst_cellmath__24_0_I734 (.Y(N1697), .A(N4149), .B(N3869));
NOR2XL inst_cellmath__24_0_I735 (.Y(N1699), .A(N4149), .B(N3877));
NOR2XL inst_cellmath__24_0_I736 (.Y(N1701), .A(N4149), .B(N3885));
NOR2XL inst_cellmath__24_0_I737 (.Y(N1703), .A(N4149), .B(N3893));
NOR2XL inst_cellmath__24_0_I738 (.Y(N1705), .A(N4149), .B(N3901));
NOR2XL inst_cellmath__24_0_I739 (.Y(N1707), .A(N4149), .B(N3909));
NOR2XL inst_cellmath__24_0_I740 (.Y(N1709), .A(N4149), .B(N3917));
NOR2XL inst_cellmath__24_0_I741 (.Y(N1711), .A(N4149), .B(N3925));
NOR2XL inst_cellmath__24_0_I742 (.Y(N1713), .A(N4149), .B(N3933));
NOR2XL inst_cellmath__24_0_I743 (.Y(N1715), .A(N4149), .B(N3941));
NOR2XL inst_cellmath__24_0_I744 (.Y(N1717), .A(N4149), .B(N3949));
NOR2XL inst_cellmath__24_0_I745 (.Y(N1719), .A(N4149), .B(N3957));
NOR2XL inst_cellmath__24_0_I746 (.Y(N1721), .A(N4149), .B(N3965));
NOR2XL inst_cellmath__24_0_I747 (.Y(N1723), .A(N4149), .B(N3973));
INVXL inst_cellmath__24_0_I748 (.Y(N1725), .A(N4149));
INVXL inst_cellmath__24_0_I754 (.Y(N1734), .A(N3793));
INVXL inst_cellmath__24_0_I755 (.Y(N1736), .A(N3805));
INVXL inst_cellmath__24_0_I756 (.Y(N1738), .A(N3813));
INVXL inst_cellmath__24_0_I757 (.Y(N1740), .A(N3820));
INVXL inst_cellmath__24_0_I758 (.Y(N1742), .A(N3826));
INVXL inst_cellmath__24_0_I759 (.Y(N1744), .A(N3834));
INVXL inst_cellmath__24_0_I760 (.Y(N1746), .A(N3845));
INVXL inst_cellmath__24_0_I761 (.Y(N1748), .A(N3853));
INVXL inst_cellmath__24_0_I762 (.Y(N1750), .A(N3861));
INVXL inst_cellmath__24_0_I763 (.Y(N1752), .A(N3869));
INVXL inst_cellmath__24_0_I764 (.Y(N1754), .A(N3877));
INVXL inst_cellmath__24_0_I765 (.Y(N1756), .A(N3885));
INVXL inst_cellmath__24_0_I766 (.Y(N1758), .A(N3893));
INVXL inst_cellmath__24_0_I767 (.Y(N1760), .A(N3901));
INVXL inst_cellmath__24_0_I768 (.Y(N1762), .A(N3909));
INVXL inst_cellmath__24_0_I769 (.Y(N1764), .A(N3917));
INVXL inst_cellmath__24_0_I770 (.Y(N1766), .A(N3925));
INVXL inst_cellmath__24_0_I771 (.Y(N1768), .A(N3933));
INVXL inst_cellmath__24_0_I772 (.Y(N1770), .A(N3941));
INVXL inst_cellmath__24_0_I773 (.Y(N1772), .A(N3949));
INVXL inst_cellmath__24_0_I774 (.Y(N1774), .A(N3957));
INVXL inst_cellmath__24_0_I775 (.Y(N1776), .A(N3965));
INVXL inst_cellmath__24_0_I776 (.Y(N1778), .A(N3973));
ADDHX1 inst_cellmath__24_0_I779 (.CO(N1783), .S(N1782), .A(N385), .B(N442));
ADDHX1 inst_cellmath__24_0_I780 (.CO(N1785), .S(N1784), .A(N387), .B(N444));
ADDFX1 inst_cellmath__24_0_I781 (.CO(N1787), .S(N1786), .A(N558), .B(N501), .CI(N1783));
ADDHX1 inst_cellmath__24_0_I782 (.CO(N1789), .S(N1788), .A(N389), .B(N446));
ADDFX1 inst_cellmath__24_0_I783 (.CO(N1791), .S(N1790), .A(N560), .B(N503), .CI(N617));
ADDFX1 inst_cellmath__24_0_I784 (.CO(N1793), .S(N1792), .A(N1788), .B(N1785), .CI(N1790));
ADDHX1 inst_cellmath__24_0_I785 (.CO(N1795), .S(N1794), .A(N391), .B(N448));
ADDFX1 inst_cellmath__24_0_I786 (.CO(N1797), .S(N1796), .A(N562), .B(N505), .CI(N619));
ADDFX1 inst_cellmath__24_0_I787 (.CO(N1799), .S(N1798), .A(N1789), .B(N676), .CI(N1794));
ADDFX1 inst_cellmath__24_0_I788 (.CO(N1801), .S(N1800), .A(N1796), .B(N1791), .CI(N1793));
ADDHX1 inst_cellmath__24_0_I789 (.CO(N1803), .S(N1802), .A(N393), .B(N450));
ADDFX1 inst_cellmath__24_0_I790 (.CO(N1805), .S(N1804), .A(N564), .B(N507), .CI(N621));
ADDFX1 inst_cellmath__24_0_I791 (.CO(N1807), .S(N1806), .A(N735), .B(N678), .CI(N1795));
ADDFX1 inst_cellmath__24_0_I792 (.CO(N1809), .S(N1808), .A(N1797), .B(N1802), .CI(N1804));
ADDFX1 inst_cellmath__24_0_I793 (.CO(N1811), .S(N1810), .A(N1806), .B(N1799), .CI(N1808));
ADDHX1 inst_cellmath__24_0_I794 (.CO(N1813), .S(N1812), .A(N395), .B(N452));
ADDFX1 inst_cellmath__24_0_I795 (.CO(N1815), .S(N1814), .A(N566), .B(N509), .CI(N623));
ADDFX1 inst_cellmath__24_0_I796 (.CO(N1817), .S(N1816), .A(N737), .B(N680), .CI(N794));
ADDFX1 inst_cellmath__24_0_I797 (.CO(N1819), .S(N1818), .A(N1812), .B(N1803), .CI(N1805));
ADDFX1 inst_cellmath__24_0_I798 (.CO(N1821), .S(N1820), .A(N1816), .B(N1814), .CI(N1807));
ADDFX1 inst_cellmath__24_0_I799 (.CO(N1823), .S(N1822), .A(N1818), .B(N1809), .CI(N1820));
ADDHX1 inst_cellmath__24_0_I800 (.CO(N1825), .S(N1824), .A(N397), .B(N454));
ADDFX1 inst_cellmath__24_0_I801 (.CO(N1827), .S(N1826), .A(N568), .B(N625), .CI(N511));
ADDFX1 inst_cellmath__24_0_I802 (.CO(N1829), .S(N1828), .A(N739), .B(N682), .CI(N796));
ADDFX1 inst_cellmath__24_0_I803 (.CO(N1831), .S(N1830), .A(N1813), .B(N853), .CI(N1824));
ADDFX1 inst_cellmath__24_0_I804 (.CO(N1833), .S(N1832), .A(N1817), .B(N1815), .CI(N1826));
ADDFX1 inst_cellmath__24_0_I805 (.CO(N1835), .S(N1834), .A(N1819), .B(N1828), .CI(N1830));
ADDFX1 inst_cellmath__24_0_I806 (.CO(N1837), .S(N1836), .A(N1832), .B(N1821), .CI(N1834));
ADDHX1 inst_cellmath__24_0_I807 (.CO(N1839), .S(N1838), .A(N399), .B(N456));
ADDFX1 inst_cellmath__24_0_I808 (.CO(N1841), .S(N1840), .A(N570), .B(N513), .CI(N627));
ADDFX1 inst_cellmath__24_0_I809 (.CO(N1843), .S(N1842), .A(N741), .B(N684), .CI(N798));
ADDFX1 inst_cellmath__24_0_I810 (.CO(N1845), .S(N1844), .A(N912), .B(N855), .CI(N1825));
ADDFX1 inst_cellmath__24_0_I811 (.CO(N1847), .S(N1846), .A(N1827), .B(N1829), .CI(N1838));
ADDFX1 inst_cellmath__24_0_I812 (.CO(N1849), .S(N1848), .A(N1842), .B(N1840), .CI(N1831));
ADDFX1 inst_cellmath__24_0_I813 (.CO(N1851), .S(N1850), .A(N1833), .B(N1844), .CI(N1846));
ADDFX1 inst_cellmath__24_0_I814 (.CO(N1853), .S(N1852), .A(N1848), .B(N1835), .CI(N1850));
ADDHX1 inst_cellmath__24_0_I815 (.CO(N1855), .S(N1854), .A(N401), .B(N458));
ADDFX1 inst_cellmath__24_0_I816 (.CO(N1857), .S(N1856), .A(N572), .B(N515), .CI(N629));
ADDFX1 inst_cellmath__24_0_I817 (.CO(N1859), .S(N1858), .A(N743), .B(N686), .CI(N800));
ADDFX1 inst_cellmath__24_0_I818 (.CO(N1861), .S(N1860), .A(N914), .B(N857), .CI(N971));
ADDFX1 inst_cellmath__24_0_I819 (.CO(N1863), .S(N1862), .A(N1854), .B(N1839), .CI(N1841));
ADDFX1 inst_cellmath__24_0_I820 (.CO(N1865), .S(N1864), .A(N1856), .B(N1843), .CI(N1845));
ADDFX1 inst_cellmath__24_0_I821 (.CO(N1867), .S(N1866), .A(N1860), .B(N1858), .CI(N1847));
ADDFX1 inst_cellmath__24_0_I822 (.CO(N1869), .S(N1868), .A(N1849), .B(N1862), .CI(N1864));
ADDFX1 inst_cellmath__24_0_I823 (.CO(N1871), .S(N1870), .A(N1851), .B(N1866), .CI(N1868));
ADDHX1 inst_cellmath__24_0_I824 (.CO(N1873), .S(N1872), .A(N403), .B(N460));
ADDFX1 inst_cellmath__24_0_I825 (.CO(N1875), .S(N1874), .A(N574), .B(N517), .CI(N631));
ADDFX1 inst_cellmath__24_0_I826 (.CO(N1877), .S(N1876), .A(N745), .B(N688), .CI(N802));
ADDFX1 inst_cellmath__24_0_I827 (.CO(N1879), .S(N1878), .A(N916), .B(N859), .CI(N973));
ADDFX1 inst_cellmath__24_0_I828 (.CO(N1881), .S(N1880), .A(N1855), .B(N1030), .CI(N1872));
ADDFX1 inst_cellmath__24_0_I829 (.CO(N1883), .S(N1882), .A(N1859), .B(N1857), .CI(N1861));
ADDFX1 inst_cellmath__24_0_I830 (.CO(N1885), .S(N1884), .A(N1876), .B(N1874), .CI(N1878));
ADDFX1 inst_cellmath__24_0_I831 (.CO(N1887), .S(N1886), .A(N1880), .B(N1863), .CI(N1882));
ADDFX1 inst_cellmath__24_0_I832 (.CO(N1889), .S(N1888), .A(N1867), .B(N1865), .CI(N1884));
ADDFX1 inst_cellmath__24_0_I833 (.CO(N1891), .S(N1890), .A(N1886), .B(N1869), .CI(N1888));
ADDHX1 inst_cellmath__24_0_I834 (.CO(N1893), .S(N1892), .A(N405), .B(N462));
ADDFX1 inst_cellmath__24_0_I835 (.CO(N1895), .S(N1894), .A(N576), .B(N519), .CI(N633));
ADDFX1 inst_cellmath__24_0_I836 (.CO(N1897), .S(N1896), .A(N747), .B(N690), .CI(N804));
ADDFX1 inst_cellmath__24_0_I837 (.CO(N1899), .S(N1898), .A(N918), .B(N861), .CI(N975));
ADDFX1 inst_cellmath__24_0_I838 (.CO(N1901), .S(N1900), .A(N1089), .B(N1032), .CI(N1873));
ADDFX1 inst_cellmath__24_0_I839 (.CO(N1903), .S(N1902), .A(N1875), .B(N1892), .CI(N1877));
ADDFX1 inst_cellmath__24_0_I840 (.CO(N1905), .S(N1904), .A(N1894), .B(N1879), .CI(N1896));
ADDFX1 inst_cellmath__24_0_I841 (.CO(N1907), .S(N1906), .A(N1881), .B(N1898), .CI(N1883));
ADDFX1 inst_cellmath__24_0_I842 (.CO(N1909), .S(N1908), .A(N1885), .B(N1900), .CI(N1902));
ADDFX1 inst_cellmath__24_0_I843 (.CO(N1911), .S(N1910), .A(N1906), .B(N1904), .CI(N1887));
ADDFX1 inst_cellmath__24_0_I844 (.CO(N1913), .S(N1912), .A(N1889), .B(N1908), .CI(N1910));
ADDHX1 inst_cellmath__24_0_I845 (.CO(N1915), .S(N1914), .A(N407), .B(N464));
ADDFX1 inst_cellmath__24_0_I846 (.CO(N1917), .S(N1916), .A(N578), .B(N521), .CI(N635));
ADDFX1 inst_cellmath__24_0_I847 (.CO(N1919), .S(N1918), .A(N749), .B(N692), .CI(N806));
ADDFX1 inst_cellmath__24_0_I848 (.CO(N1921), .S(N1920), .A(N920), .B(N863), .CI(N977));
ADDFX1 inst_cellmath__24_0_I849 (.CO(N1923), .S(N1922), .A(N1091), .B(N1034), .CI(N1148));
ADDFX1 inst_cellmath__24_0_I850 (.CO(N1925), .S(N1924), .A(N1914), .B(N1893), .CI(N1895));
ADDFX1 inst_cellmath__24_0_I851 (.CO(N1927), .S(N1926), .A(N1899), .B(N1897), .CI(N1916));
ADDFX1 inst_cellmath__24_0_I852 (.CO(N1929), .S(N1928), .A(N1920), .B(N1918), .CI(N1901));
ADDFX1 inst_cellmath__24_0_I853 (.CO(N1931), .S(N1930), .A(N1903), .B(N1922), .CI(N1905));
ADDFX1 inst_cellmath__24_0_I854 (.CO(N1933), .S(N1932), .A(N1926), .B(N1924), .CI(N1928));
ADDFX1 inst_cellmath__24_0_I855 (.CO(N1935), .S(N1934), .A(N1909), .B(N1907), .CI(N1930));
ADDFX1 inst_cellmath__24_0_I856 (.CO(N1937), .S(N1936), .A(N1911), .B(N1932), .CI(N1934));
ADDHX1 inst_cellmath__24_0_I857 (.CO(N1939), .S(N1938), .A(N409), .B(N466));
ADDFX1 inst_cellmath__24_0_I858 (.CO(N1941), .S(N1940), .A(N580), .B(N523), .CI(N637));
ADDFX1 inst_cellmath__24_0_I859 (.CO(N1943), .S(N1942), .A(N751), .B(N694), .CI(N808));
ADDFX1 inst_cellmath__24_0_I860 (.CO(N1945), .S(N1944), .A(N922), .B(N865), .CI(N979));
ADDFX1 inst_cellmath__24_0_I861 (.CO(N1947), .S(N1946), .A(N1093), .B(N1036), .CI(N1150));
ADDFX1 inst_cellmath__24_0_I862 (.CO(N1949), .S(N1948), .A(N1915), .B(N1207), .CI(N1938));
ADDFX1 inst_cellmath__24_0_I863 (.CO(N1951), .S(N1950), .A(N1919), .B(N1917), .CI(N1921));
ADDFX1 inst_cellmath__24_0_I864 (.CO(N1953), .S(N1952), .A(N1940), .B(N1923), .CI(N1942));
ADDFX1 inst_cellmath__24_0_I865 (.CO(N1955), .S(N1954), .A(N1946), .B(N1944), .CI(N1925));
ADDFX1 inst_cellmath__24_0_I866 (.CO(N1957), .S(N1956), .A(N1948), .B(N1927), .CI(N1950));
ADDFX1 inst_cellmath__24_0_I867 (.CO(N1959), .S(N1958), .A(N1952), .B(N1929), .CI(N1931));
ADDFXL inst_cellmath__24_0_I868 (.CO(N1961), .S(N1960), .A(N1933), .B(N1954), .CI(N1956));
ADDFX1 inst_cellmath__24_0_I869 (.CO(N1963), .S(N1962), .A(N1958), .B(N1935), .CI(N1960));
ADDHX1 inst_cellmath__24_0_I870 (.CO(N1965), .S(N1964), .A(N411), .B(N468));
ADDFX1 inst_cellmath__24_0_I871 (.CO(N1967), .S(N1966), .A(N582), .B(N525), .CI(N639));
ADDFX1 inst_cellmath__24_0_I872 (.CO(N1969), .S(N1968), .A(N753), .B(N696), .CI(N810));
ADDFX1 inst_cellmath__24_0_I873 (.CO(N1971), .S(N1970), .A(N924), .B(N867), .CI(N981));
ADDFX1 inst_cellmath__24_0_I874 (.CO(N1973), .S(N1972), .A(N1095), .B(N1038), .CI(N1152));
ADDFX1 inst_cellmath__24_0_I875 (.CO(N1975), .S(N1974), .A(N1266), .B(N1209), .CI(N1939));
ADDFX1 inst_cellmath__24_0_I876 (.CO(N1977), .S(N1976), .A(N1941), .B(N1964), .CI(N1943));
ADDFX1 inst_cellmath__24_0_I877 (.CO(N1979), .S(N1978), .A(N1947), .B(N1945), .CI(N1966));
ADDFX1 inst_cellmath__24_0_I878 (.CO(N1981), .S(N1980), .A(N1970), .B(N1968), .CI(N1972));
ADDFX1 inst_cellmath__24_0_I879 (.CO(N1983), .S(N1982), .A(N1974), .B(N1949), .CI(N1951));
ADDFX1 inst_cellmath__24_0_I880 (.CO(N1985), .S(N1984), .A(N1976), .B(N1953), .CI(N1978));
ADDFX1 inst_cellmath__24_0_I881 (.CO(N1987), .S(N1986), .A(N1955), .B(N1980), .CI(N1982));
ADDFX1 inst_cellmath__24_0_I882 (.CO(N1989), .S(N1988), .A(N1984), .B(N1957), .CI(N1959));
ADDFX1 inst_cellmath__24_0_I883 (.CO(N1991), .S(N1990), .A(N1961), .B(N1986), .CI(N1988));
ADDHX1 inst_cellmath__24_0_I884 (.CO(N1993), .S(N1992), .A(N413), .B(N470));
ADDFX1 inst_cellmath__24_0_I885 (.CO(N1995), .S(N1994), .A(N584), .B(N527), .CI(N641));
ADDFX1 inst_cellmath__24_0_I886 (.CO(N1997), .S(N1996), .A(N755), .B(N698), .CI(N812));
ADDFX1 inst_cellmath__24_0_I887 (.CO(N1999), .S(N1998), .A(N926), .B(N869), .CI(N983));
ADDFX1 inst_cellmath__24_0_I888 (.CO(N2001), .S(N2000), .A(N1097), .B(N1040), .CI(N1154));
ADDFX1 inst_cellmath__24_0_I889 (.CO(N2003), .S(N2002), .A(N1268), .B(N1211), .CI(N1325));
ADDFX1 inst_cellmath__24_0_I890 (.CO(N2005), .S(N2004), .A(N1992), .B(N1965), .CI(N1967));
ADDFX1 inst_cellmath__24_0_I891 (.CO(N2007), .S(N2006), .A(N1971), .B(N1969), .CI(N1973));
ADDFX1 inst_cellmath__24_0_I892 (.CO(N2009), .S(N2008), .A(N1996), .B(N1994), .CI(N1975));
ADDFX1 inst_cellmath__24_0_I893 (.CO(N2011), .S(N2010), .A(N2000), .B(N1998), .CI(N2002));
ADDFX1 inst_cellmath__24_0_I894 (.CO(N2013), .S(N2012), .A(N1979), .B(N1977), .CI(N1981));
ADDFX1 inst_cellmath__24_0_I895 (.CO(N2015), .S(N2014), .A(N2004), .B(N2006), .CI(N2008));
ADDFX1 inst_cellmath__24_0_I896 (.CO(N2017), .S(N2016), .A(N1983), .B(N2010), .CI(N1985));
ADDFX1 inst_cellmath__24_0_I897 (.CO(N2019), .S(N2018), .A(N2014), .B(N2012), .CI(N1987));
ADDFX1 inst_cellmath__24_0_I898 (.CO(N2021), .S(N2020), .A(N1989), .B(N2016), .CI(N2018));
ADDHX1 inst_cellmath__24_0_I899 (.CO(N2023), .S(N2022), .A(N415), .B(N472));
ADDFX1 inst_cellmath__24_0_I900 (.CO(N2025), .S(N2024), .A(N643), .B(N529), .CI(N586));
ADDFX1 inst_cellmath__24_0_I901 (.CO(N2027), .S(N2026), .A(N757), .B(N700), .CI(N814));
ADDFX1 inst_cellmath__24_0_I902 (.CO(N2029), .S(N2028), .A(N928), .B(N871), .CI(N985));
ADDFX1 inst_cellmath__24_0_I903 (.CO(N2031), .S(N2030), .A(N1099), .B(N1042), .CI(N1156));
ADDFX1 inst_cellmath__24_0_I904 (.CO(N2033), .S(N2032), .A(N1270), .B(N1213), .CI(N1327));
ADDFX1 inst_cellmath__24_0_I905 (.CO(N2035), .S(N2034), .A(N1993), .B(N1384), .CI(N2022));
ADDFX1 inst_cellmath__24_0_I906 (.CO(N2037), .S(N2036), .A(N1997), .B(N1995), .CI(N1999));
ADDFX1 inst_cellmath__24_0_I907 (.CO(N2039), .S(N2038), .A(N2001), .B(N2003), .CI(N2024));
ADDFXL inst_cellmath__24_0_I908 (.CO(N2041), .S(N2040), .A(N2028), .B(N2026), .CI(N2030));
ADDFX1 inst_cellmath__24_0_I909 (.CO(N2043), .S(N2042), .A(N2007), .B(N2032), .CI(N2005));
ADDFX1 inst_cellmath__24_0_I910 (.CO(N2045), .S(N2044), .A(N2009), .B(N2034), .CI(N2036));
ADDFX1 inst_cellmath__24_0_I911 (.CO(N2047), .S(N2046), .A(N2038), .B(N2011), .CI(N2040));
ADDFX1 inst_cellmath__24_0_I912 (.CO(N2049), .S(N2048), .A(N2042), .B(N2013), .CI(N2015));
ADDFHXL inst_cellmath__24_0_I913 (.CO(N2051), .S(N2050), .A(N2046), .B(N2044), .CI(N2017));
ADDFHXL inst_cellmath__24_0_I914 (.CO(N2053), .S(N2052), .A(N2019), .B(N2048), .CI(N2050));
ADDHX1 inst_cellmath__24_0_I915 (.CO(N2055), .S(N2054), .A(N417), .B(N474));
ADDFX1 inst_cellmath__24_0_I916 (.CO(N2057), .S(N2056), .A(N588), .B(N531), .CI(N645));
ADDFX1 inst_cellmath__24_0_I917 (.CO(N2059), .S(N2058), .A(N759), .B(N702), .CI(N816));
ADDFX1 inst_cellmath__24_0_I918 (.CO(N2061), .S(N2060), .A(N930), .B(N873), .CI(N987));
ADDFX1 inst_cellmath__24_0_I919 (.CO(N2063), .S(N2062), .A(N1101), .B(N1044), .CI(N1158));
ADDFX1 inst_cellmath__24_0_I920 (.CO(N2065), .S(N2064), .A(N1272), .B(N1215), .CI(N1329));
ADDFX1 inst_cellmath__24_0_I921 (.CO(N2067), .S(N2066), .A(N1443), .B(N1386), .CI(N2023));
ADDFX1 inst_cellmath__24_0_I922 (.CO(N2069), .S(N2068), .A(N2025), .B(N2054), .CI(N2027));
ADDFX1 inst_cellmath__24_0_I923 (.CO(N2071), .S(N2070), .A(N2031), .B(N2029), .CI(N2033));
ADDFX1 inst_cellmath__24_0_I924 (.CO(N2073), .S(N2072), .A(N2058), .B(N2056), .CI(N2060));
ADDFX1 inst_cellmath__24_0_I925 (.CO(N2075), .S(N2074), .A(N2064), .B(N2062), .CI(N2035));
ADDFX1 inst_cellmath__24_0_I926 (.CO(N2077), .S(N2076), .A(N2037), .B(N2066), .CI(N2039));
ADDFX1 inst_cellmath__24_0_I927 (.CO(N2079), .S(N2078), .A(N2070), .B(N2041), .CI(N2068));
ADDFX1 inst_cellmath__24_0_I928 (.CO(N2081), .S(N2080), .A(N2043), .B(N2072), .CI(N2074));
ADDFX1 inst_cellmath__24_0_I929 (.CO(N2083), .S(N2082), .A(N2076), .B(N2045), .CI(N2047));
ADDFX1 inst_cellmath__24_0_I930 (.CO(N2085), .S(N2084), .A(N2080), .B(N2078), .CI(N2049));
ADDFHXL inst_cellmath__24_0_I931 (.CO(N2087), .S(N2086), .A(N2051), .B(N2082), .CI(N2084));
ADDHX1 inst_cellmath__24_0_I932 (.CO(N2089), .S(N2088), .A(N419), .B(N476));
ADDFX1 inst_cellmath__24_0_I933 (.CO(N2091), .S(N2090), .A(N590), .B(N533), .CI(N647));
ADDFX1 inst_cellmath__24_0_I934 (.CO(N2093), .S(N2092), .A(N761), .B(N704), .CI(N818));
ADDFX1 inst_cellmath__24_0_I935 (.CO(N2095), .S(N2094), .A(N932), .B(N875), .CI(N989));
ADDFX1 inst_cellmath__24_0_I936 (.CO(N2097), .S(N2096), .A(N1103), .B(N1046), .CI(N1160));
ADDFX1 inst_cellmath__24_0_I937 (.CO(N2099), .S(N2098), .A(N1274), .B(N1217), .CI(N1331));
ADDFX1 inst_cellmath__24_0_I938 (.CO(N2101), .S(N2100), .A(N1445), .B(N1388), .CI(N1502));
ADDFX1 inst_cellmath__24_0_I939 (.CO(N2103), .S(N2102), .A(N2088), .B(N2055), .CI(N2057));
ADDFX1 inst_cellmath__24_0_I940 (.CO(N2105), .S(N2104), .A(N2061), .B(N2059), .CI(N2063));
ADDFX1 inst_cellmath__24_0_I941 (.CO(N2107), .S(N2106), .A(N2090), .B(N2065), .CI(N2067));
ADDFX1 inst_cellmath__24_0_I942 (.CO(N2109), .S(N2108), .A(N2094), .B(N2092), .CI(N2096));
ADDFXL inst_cellmath__24_0_I943 (.CO(N2111), .S(N2110), .A(N2100), .B(N2098), .CI(N2069));
ADDFX1 inst_cellmath__24_0_I944 (.CO(N2113), .S(N2112), .A(N2073), .B(N2071), .CI(N2102));
ADDFX1 inst_cellmath__24_0_I945 (.CO(N2115), .S(N2114), .A(N2075), .B(N2104), .CI(N2106));
ADDFXL inst_cellmath__24_0_I946 (.CO(N2117), .S(N2116), .A(N2077), .B(N2108), .CI(N2110));
ADDFX1 inst_cellmath__24_0_I947 (.CO(N2119), .S(N2118), .A(N2112), .B(N2079), .CI(N2081));
ADDFXL inst_cellmath__24_0_I948 (.CO(N2121), .S(N2120), .A(N2116), .B(N2114), .CI(N2083));
ADDFX1 inst_cellmath__24_0_I949 (.CO(N2123), .S(N2122), .A(N2085), .B(N2118), .CI(N2120));
ADDHX1 inst_cellmath__24_0_I950 (.CO(N2125), .S(N2124), .A(N421), .B(N478));
ADDFX1 inst_cellmath__24_0_I951 (.CO(N2127), .S(N2126), .A(N592), .B(N535), .CI(N649));
ADDFX1 inst_cellmath__24_0_I952 (.CO(N2129), .S(N2128), .A(N763), .B(N706), .CI(N820));
ADDFXL inst_cellmath__24_0_I953 (.CO(N2131), .S(N2130), .A(N934), .B(N877), .CI(N991));
ADDFX1 inst_cellmath__24_0_I954 (.CO(N2133), .S(N2132), .A(N1105), .B(N1048), .CI(N1162));
ADDFX1 inst_cellmath__24_0_I955 (.CO(N2135), .S(N2134), .A(N1276), .B(N1219), .CI(N1333));
ADDFX1 inst_cellmath__24_0_I956 (.CO(N2137), .S(N2136), .A(N1447), .B(N1390), .CI(N1504));
ADDFX1 inst_cellmath__24_0_I957 (.CO(N2139), .S(N2138), .A(N2089), .B(N1561), .CI(N2124));
ADDFX1 inst_cellmath__24_0_I958 (.CO(N2141), .S(N2140), .A(N2093), .B(N2091), .CI(N2095));
ADDFX1 inst_cellmath__24_0_I959 (.CO(N2143), .S(N2142), .A(N2099), .B(N2097), .CI(N2101));
ADDFX1 inst_cellmath__24_0_I960 (.CO(N2145), .S(N2144), .A(N2128), .B(N2126), .CI(N2130));
ADDFX1 inst_cellmath__24_0_I961 (.CO(N2147), .S(N2146), .A(N2134), .B(N2132), .CI(N2136));
ADDFX1 inst_cellmath__24_0_I962 (.CO(N2149), .S(N2148), .A(N2103), .B(N2105), .CI(N2138));
ADDFX1 inst_cellmath__24_0_I963 (.CO(N2151), .S(N2150), .A(N2140), .B(N2142), .CI(N2107));
ADDFX1 inst_cellmath__24_0_I964 (.CO(N2153), .S(N2152), .A(N2111), .B(N2109), .CI(N2144));
ADDFX1 inst_cellmath__24_0_I965 (.CO(N2155), .S(N2154), .A(N2113), .B(N2146), .CI(N2148));
ADDFX1 inst_cellmath__24_0_I966 (.CO(N2157), .S(N2156), .A(N2150), .B(N2115), .CI(N2117));
ADDFX1 inst_cellmath__24_0_I967 (.CO(N2159), .S(N2158), .A(N2154), .B(N2152), .CI(N2119));
ADDFXL inst_cellmath__24_0_I968 (.CO(N2161), .S(N2160), .A(N2121), .B(N2156), .CI(N2158));
ADDHX1 inst_cellmath__24_0_I969 (.CO(N2163), .S(N2162), .A(N423), .B(N480));
ADDFX1 inst_cellmath__24_0_I970 (.CO(N2165), .S(N2164), .A(N594), .B(N537), .CI(N651));
ADDFX1 inst_cellmath__24_0_I971 (.CO(N2167), .S(N2166), .A(N822), .B(N708), .CI(N765));
ADDFX1 inst_cellmath__24_0_I972 (.CO(N2169), .S(N2168), .A(N936), .B(N879), .CI(N993));
ADDFX1 inst_cellmath__24_0_I973 (.CO(N2171), .S(N2170), .A(N1107), .B(N1050), .CI(N1164));
ADDFX1 inst_cellmath__24_0_I974 (.CO(N2173), .S(N2172), .A(N1278), .B(N1221), .CI(N1335));
ADDFX1 inst_cellmath__24_0_I975 (.CO(N2175), .S(N2174), .A(N1449), .B(N1392), .CI(N1506));
ADDFX1 inst_cellmath__24_0_I976 (.CO(N2177), .S(N2176), .A(N1563), .B(N1620), .CI(N2125));
ADDFX1 inst_cellmath__24_0_I977 (.CO(N2179), .S(N2178), .A(N2127), .B(N2162), .CI(N2129));
ADDFX1 inst_cellmath__24_0_I978 (.CO(N2181), .S(N2180), .A(N2133), .B(N2131), .CI(N2135));
ADDFX1 inst_cellmath__24_0_I979 (.CO(N2183), .S(N2182), .A(N2164), .B(N2137), .CI(N2166));
ADDFX1 inst_cellmath__24_0_I980 (.CO(N2185), .S(N2184), .A(N2170), .B(N2168), .CI(N2172));
ADDFX1 inst_cellmath__24_0_I981 (.CO(N2187), .S(N2186), .A(N2139), .B(N2174), .CI(N2141));
ADDFHXL inst_cellmath__24_0_I982 (.CO(N2189), .S(N2188), .A(N2143), .B(N2176), .CI(N2145));
ADDFX1 inst_cellmath__24_0_I983 (.CO(N2191), .S(N2190), .A(N2180), .B(N2147), .CI(N2178));
ADDFXL inst_cellmath__24_0_I984 (.CO(N2193), .S(N2192), .A(N2184), .B(N2182), .CI(N2149));
ADDFHXL inst_cellmath__24_0_I985 (.CO(N2195), .S(N2194), .A(N2151), .B(N2186), .CI(N2188));
ADDFX1 inst_cellmath__24_0_I986 (.CO(N2197), .S(N2196), .A(N2190), .B(N2153), .CI(N2192));
ADDFX1 inst_cellmath__24_0_I987 (.CO(N2199), .S(N2198), .A(N2194), .B(N2155), .CI(N2157));
ADDFXL inst_cellmath__24_0_I988 (.CO(N2201), .S(N2200), .A(N2159), .B(N2196), .CI(N2198));
ADDHX1 inst_cellmath__24_0_I989 (.CO(N2203), .S(N2202), .A(N425), .B(N482));
ADDFXL inst_cellmath__24_0_I990 (.CO(N2205), .S(N2204), .A(N653), .B(N539), .CI(N596));
ADDFX1 inst_cellmath__24_0_I991 (.CO(N2207), .S(N2206), .A(N824), .B(N710), .CI(N767));
ADDFX1 inst_cellmath__24_0_I992 (.CO(N2209), .S(N2208), .A(N995), .B(N938), .CI(N881));
ADDFX1 inst_cellmath__24_0_I993 (.CO(N2211), .S(N2210), .A(N1109), .B(N1052), .CI(N1166));
ADDFX1 inst_cellmath__24_0_I994 (.CO(N2213), .S(N2212), .A(N1280), .B(N1337), .CI(N1223));
ADDFX1 inst_cellmath__24_0_I995 (.CO(N2215), .S(N2214), .A(N1451), .B(N1508), .CI(N1394));
ADDFX1 inst_cellmath__24_0_I996 (.CO(N2217), .S(N2216), .A(N1622), .B(N1565), .CI(N1679));
ADDFX1 inst_cellmath__24_0_I997 (.CO(N2219), .S(N2218), .A(N2202), .B(N2163), .CI(N2165));
ADDFX1 inst_cellmath__24_0_I998 (.CO(N2221), .S(N2220), .A(N2169), .B(N2167), .CI(N2171));
ADDFXL inst_cellmath__24_0_I999 (.CO(N2223), .S(N2222), .A(N2175), .B(N2173), .CI(N2204));
ADDFHXL inst_cellmath__24_0_I1000 (.CO(N2225), .S(N2224), .A(N2208), .B(N2206), .CI(N2177));
ADDFX1 inst_cellmath__24_0_I1001 (.CO(N2227), .S(N2226), .A(N2212), .B(N2210), .CI(N2214));
ADDFX1 inst_cellmath__24_0_I1002 (.CO(N2229), .S(N2228), .A(N2179), .B(N2216), .CI(N2181));
ADDFXL inst_cellmath__24_0_I1003 (.CO(N2231), .S(N2230), .A(N2220), .B(N2218), .CI(N2183));
ADDFX1 inst_cellmath__24_0_I1004 (.CO(N2233), .S(N2232), .A(N2222), .B(N2185), .CI(N2224));
ADDFX1 inst_cellmath__24_0_I1005 (.CO(N2235), .S(N2234), .A(N2226), .B(N2187), .CI(N2189));
ADDFX1 inst_cellmath__24_0_I1006 (.CO(N2237), .S(N2236), .A(N2228), .B(N2191), .CI(N2230));
ADDFHXL inst_cellmath__24_0_I1007 (.CO(N2239), .S(N2238), .A(N2232), .B(N2193), .CI(N2195));
ADDFHXL inst_cellmath__24_0_I1008 (.CO(N2241), .S(N2240), .A(N2236), .B(N2234), .CI(N2197));
ADDFHXL inst_cellmath__24_0_I1009 (.CO(N2243), .S(N2242), .A(N2199), .B(N2238), .CI(N2240));
ADDHX1 inst_cellmath__24_0_I1010 (.CO(N2245), .S(N2244), .A(N1734), .B(N484));
ADDFX1 inst_cellmath__24_0_I1011 (.CO(N2247), .S(N2246), .A(N541), .B(N427), .CI(N598));
ADDFX1 inst_cellmath__24_0_I1012 (.CO(N2249), .S(N2248), .A(N712), .B(N655), .CI(N769));
ADDFX1 inst_cellmath__24_0_I1013 (.CO(N2251), .S(N2250), .A(N883), .B(N826), .CI(N940));
ADDFX1 inst_cellmath__24_0_I1014 (.CO(N2253), .S(N2252), .A(N1054), .B(N997), .CI(N1111));
ADDFX1 inst_cellmath__24_0_I1015 (.CO(N2255), .S(N2254), .A(N1225), .B(N1168), .CI(N1282));
ADDFX1 inst_cellmath__24_0_I1016 (.CO(N2257), .S(N2256), .A(N1396), .B(N1339), .CI(N1453));
ADDFX1 inst_cellmath__24_0_I1017 (.CO(N2259), .S(N2258), .A(N1567), .B(N1510), .CI(N1624));
ADDFHXL inst_cellmath__24_0_I1018 (.CO(N2261), .S(N2260), .A(N2203), .B(N1681), .CI(N2244));
ADDFX1 inst_cellmath__24_0_I1019 (.CO(N2263), .S(N2262), .A(N2209), .B(N2205), .CI(N2207));
ADDFXL inst_cellmath__24_0_I1020 (.CO(N2265), .S(N2264), .A(N2213), .B(N2215), .CI(N2211));
ADDFX1 inst_cellmath__24_0_I1021 (.CO(N2267), .S(N2266), .A(N2246), .B(N2217), .CI(N2248));
ADDFX1 inst_cellmath__24_0_I1022 (.CO(N2269), .S(N2268), .A(N2252), .B(N2250), .CI(N2254));
ADDFXL inst_cellmath__24_0_I1023 (.CO(N2271), .S(N2270), .A(N2258), .B(N2256), .CI(N2221));
ADDFX1 inst_cellmath__24_0_I1024 (.CO(N2273), .S(N2272), .A(N2260), .B(N2219), .CI(N2223));
ADDFXL inst_cellmath__24_0_I1025 (.CO(N2275), .S(N2274), .A(N2225), .B(N2262), .CI(N2264));
ADDFX1 inst_cellmath__24_0_I1026 (.CO(N2277), .S(N2276), .A(N2266), .B(N2227), .CI(N2268));
ADDFXL inst_cellmath__24_0_I1027 (.CO(N2279), .S(N2278), .A(N2270), .B(N2229), .CI(N2231));
ADDFHXL inst_cellmath__24_0_I1028 (.CO(N2281), .S(N2280), .A(N2233), .B(N2272), .CI(N2274));
ADDFX1 inst_cellmath__24_0_I1029 (.CO(N2283), .S(N2282), .A(N2276), .B(N2235), .CI(N2278));
ADDFHXL inst_cellmath__24_0_I1030 (.CO(N2285), .S(N2284), .A(N2280), .B(N2237), .CI(N2239));
ADDFHX1 inst_cellmath__24_0_I1031 (.CO(N2287), .S(N2286), .A(N2241), .B(N2282), .CI(N2284));
ADDHX1 inst_cellmath__24_0_I1032 (.CO(N2289), .S(N2288), .A(N1736), .B(N543));
ADDFXL inst_cellmath__24_0_I1033 (.CO(N2291), .S(N2290), .A(N657), .B(N486), .CI(N600));
ADDFX1 inst_cellmath__24_0_I1034 (.CO(N2293), .S(N2292), .A(N714), .B(N771), .CI(N828));
ADDFX1 inst_cellmath__24_0_I1035 (.CO(N2295), .S(N2294), .A(N942), .B(N885), .CI(N999));
ADDFX1 inst_cellmath__24_0_I1036 (.CO(N2297), .S(N2296), .A(N1113), .B(N1056), .CI(N1170));
ADDFX1 inst_cellmath__24_0_I1037 (.CO(N2299), .S(N2298), .A(N1284), .B(N1227), .CI(N1341));
ADDFX1 inst_cellmath__24_0_I1038 (.CO(N2301), .S(N2300), .A(N1455), .B(N1398), .CI(N1512));
ADDFX1 inst_cellmath__24_0_I1039 (.CO(N2303), .S(N2302), .A(N1626), .B(N1569), .CI(N1683));
ADDFX1 inst_cellmath__24_0_I1040 (.CO(N2305), .S(N2304), .A(N2288), .B(N2245), .CI(N2247));
ADDFX1 inst_cellmath__24_0_I1041 (.CO(N2307), .S(N2306), .A(N2251), .B(N2249), .CI(N2253));
ADDFX1 inst_cellmath__24_0_I1042 (.CO(N2309), .S(N2308), .A(N2257), .B(N2255), .CI(N2259));
ADDFXL inst_cellmath__24_0_I1043 (.CO(N2311), .S(N2310), .A(N2292), .B(N2290), .CI(N2294));
ADDFX1 inst_cellmath__24_0_I1044 (.CO(N2313), .S(N2312), .A(N2298), .B(N2296), .CI(N2300));
ADDFHXL inst_cellmath__24_0_I1045 (.CO(N2315), .S(N2314), .A(N2261), .B(N2302), .CI(N2263));
ADDFX1 inst_cellmath__24_0_I1046 (.CO(N2317), .S(N2316), .A(N2304), .B(N2265), .CI(N2306));
ADDFXL inst_cellmath__24_0_I1047 (.CO(N2319), .S(N2318), .A(N2308), .B(N2267), .CI(N2269));
ADDFX1 inst_cellmath__24_0_I1048 (.CO(N2321), .S(N2320), .A(N2310), .B(N2271), .CI(N2312));
ADDFHXL inst_cellmath__24_0_I1049 (.CO(N2323), .S(N2322), .A(N2273), .B(N2314), .CI(N2275));
ADDFHXL inst_cellmath__24_0_I1050 (.CO(N2325), .S(N2324), .A(N2318), .B(N2316), .CI(N2277));
ADDFHXL inst_cellmath__24_0_I1051 (.CO(N2327), .S(N2326), .A(N2320), .B(N2279), .CI(N2322));
ADDFHXL inst_cellmath__24_0_I1052 (.CO(N2329), .S(N2328), .A(N2324), .B(N2281), .CI(N2283));
ADDFHXL inst_cellmath__24_0_I1053 (.CO(N2331), .S(N2330), .A(N2285), .B(N2326), .CI(N2328));
ADDFX1 inst_cellmath__24_0_I1054 (.CO(N2333), .S(N2332), .A(N545), .B(N1738), .CI(N602));
ADDFX1 inst_cellmath__24_0_I1055 (.CO(N2335), .S(N2334), .A(N716), .B(N659), .CI(N773));
ADDFX1 inst_cellmath__24_0_I1056 (.CO(N2337), .S(N2336), .A(N887), .B(N830), .CI(N944));
ADDFX1 inst_cellmath__24_0_I1057 (.CO(N2339), .S(N2338), .A(N1058), .B(N1001), .CI(N1115));
ADDFX1 inst_cellmath__24_0_I1058 (.CO(N2341), .S(N2340), .A(N1229), .B(N1172), .CI(N1286));
ADDFX1 inst_cellmath__24_0_I1059 (.CO(N2343), .S(N2342), .A(N1400), .B(N1343), .CI(N1457));
ADDFX1 inst_cellmath__24_0_I1060 (.CO(N2345), .S(N2344), .A(N1571), .B(N1514), .CI(N1628));
ADDFXL inst_cellmath__24_0_I1061 (.CO(N2347), .S(N2346), .A(N2289), .B(N1685), .CI(N2291));
ADDFX1 inst_cellmath__24_0_I1062 (.CO(N2349), .S(N2348), .A(N2295), .B(N2293), .CI(N2297));
ADDFX1 inst_cellmath__24_0_I1063 (.CO(N2351), .S(N2350), .A(N2301), .B(N2299), .CI(N2303));
ADDFX1 inst_cellmath__24_0_I1064 (.CO(N2353), .S(N2352), .A(N2334), .B(N2332), .CI(N2336));
ADDFX1 inst_cellmath__24_0_I1065 (.CO(N2355), .S(N2354), .A(N2340), .B(N2338), .CI(N2342));
ADDFHXL inst_cellmath__24_0_I1066 (.CO(N2357), .S(N2356), .A(N2305), .B(N2344), .CI(N2307));
ADDFX1 inst_cellmath__24_0_I1067 (.CO(N2359), .S(N2358), .A(N2346), .B(N2309), .CI(N2311));
ADDFXL inst_cellmath__24_0_I1068 (.CO(N2361), .S(N2360), .A(N2348), .B(N2313), .CI(N2350));
ADDFX1 inst_cellmath__24_0_I1069 (.CO(N2363), .S(N2362), .A(N2354), .B(N2315), .CI(N2352));
ADDFHXL inst_cellmath__24_0_I1070 (.CO(N2365), .S(N2364), .A(N2356), .B(N2317), .CI(N2319));
ADDFHXL inst_cellmath__24_0_I1071 (.CO(N2367), .S(N2366), .A(N2360), .B(N2358), .CI(N2321));
ADDFXL inst_cellmath__24_0_I1072 (.CO(N2369), .S(N2368), .A(N2362), .B(N2323), .CI(N2364));
ADDFHXL inst_cellmath__24_0_I1073 (.CO(N2371), .S(N2370), .A(N2366), .B(N2325), .CI(N2327));
ADDFHXL inst_cellmath__24_0_I1074 (.CO(N2373), .S(N2372), .A(N2329), .B(N2368), .CI(N2370));
ADDFX1 inst_cellmath__24_0_I1075 (.CO(N2375), .S(N2374), .A(N604), .B(N1740), .CI(N661));
ADDFX1 inst_cellmath__24_0_I1076 (.CO(N2377), .S(N2376), .A(N775), .B(N718), .CI(N832));
ADDFX1 inst_cellmath__24_0_I1077 (.CO(N2379), .S(N2378), .A(N946), .B(N889), .CI(N1003));
ADDFX1 inst_cellmath__24_0_I1078 (.CO(N2381), .S(N2380), .A(N1117), .B(N1060), .CI(N1174));
ADDFX1 inst_cellmath__24_0_I1079 (.CO(N2383), .S(N2382), .A(N1288), .B(N1231), .CI(N1345));
ADDFX1 inst_cellmath__24_0_I1080 (.CO(N2385), .S(N2384), .A(N1459), .B(N1402), .CI(N1516));
ADDFX1 inst_cellmath__24_0_I1081 (.CO(N2387), .S(N2386), .A(N1630), .B(N1573), .CI(N1687));
ADDFX1 inst_cellmath__24_0_I1082 (.CO(N2389), .S(N2388), .A(N2335), .B(N2333), .CI(N2337));
ADDFX1 inst_cellmath__24_0_I1083 (.CO(N2391), .S(N2390), .A(N2341), .B(N2339), .CI(N2343));
ADDFX1 inst_cellmath__24_0_I1084 (.CO(N2393), .S(N2392), .A(N2374), .B(N2345), .CI(N2376));
ADDFXL inst_cellmath__24_0_I1085 (.CO(N2395), .S(N2394), .A(N2380), .B(N2378), .CI(N2382));
ADDFX1 inst_cellmath__24_0_I1086 (.CO(N2397), .S(N2396), .A(N2386), .B(N2384), .CI(N2347));
ADDFHX1 inst_cellmath__24_0_I1087 (.CO(N2399), .S(N2398), .A(N2351), .B(N2349), .CI(N2353));
ADDFXL inst_cellmath__24_0_I1088 (.CO(N2401), .S(N2400), .A(N2388), .B(N2355), .CI(N2390));
ADDFHXL inst_cellmath__24_0_I1089 (.CO(N2403), .S(N2402), .A(N2394), .B(N2392), .CI(N2357));
ADDFHXL inst_cellmath__24_0_I1090 (.CO(N2405), .S(N2404), .A(N2359), .B(N2396), .CI(N2361));
ADDFX1 inst_cellmath__24_0_I1091 (.CO(N2407), .S(N2406), .A(N2400), .B(N2398), .CI(N2363));
ADDFHXL inst_cellmath__24_0_I1092 (.CO(N2409), .S(N2408), .A(N2402), .B(N2365), .CI(N2404));
ADDFHXL inst_cellmath__24_0_I1093 (.CO(N2411), .S(N2410), .A(N2406), .B(N2367), .CI(N2369));
ADDFHXL inst_cellmath__24_0_I1094 (.CO(N2413), .S(N2412), .A(N2371), .B(N2408), .CI(N2410));
ADDFX1 inst_cellmath__24_0_I1095 (.CO(N2415), .S(N2414), .A(N663), .B(N1742), .CI(N720));
ADDFX1 inst_cellmath__24_0_I1096 (.CO(N2417), .S(N2416), .A(N834), .B(N777), .CI(N891));
ADDFX1 inst_cellmath__24_0_I1097 (.CO(N2419), .S(N2418), .A(N1005), .B(N948), .CI(N1062));
ADDFX1 inst_cellmath__24_0_I1098 (.CO(N2421), .S(N2420), .A(N1176), .B(N1119), .CI(N1233));
ADDFX1 inst_cellmath__24_0_I1099 (.CO(N2423), .S(N2422), .A(N1347), .B(N1290), .CI(N1404));
ADDFX1 inst_cellmath__24_0_I1100 (.CO(N2425), .S(N2424), .A(N1518), .B(N1461), .CI(N1575));
ADDFX1 inst_cellmath__24_0_I1101 (.CO(N2427), .S(N2426), .A(N1689), .B(N1632), .CI(N2375));
ADDFX1 inst_cellmath__24_0_I1102 (.CO(N2429), .S(N2428), .A(N2379), .B(N2377), .CI(N2381));
ADDFX1 inst_cellmath__24_0_I1103 (.CO(N2431), .S(N2430), .A(N2385), .B(N2383), .CI(N2387));
ADDFX1 inst_cellmath__24_0_I1104 (.CO(N2433), .S(N2432), .A(N2416), .B(N2414), .CI(N2418));
ADDFX1 inst_cellmath__24_0_I1105 (.CO(N2435), .S(N2434), .A(N2422), .B(N2420), .CI(N2424));
ADDFX1 inst_cellmath__24_0_I1106 (.CO(N2437), .S(N2436), .A(N2391), .B(N2389), .CI(N2426));
ADDFHXL inst_cellmath__24_0_I1107 (.CO(N2439), .S(N2438), .A(N2428), .B(N2393), .CI(N2395));
ADDFX1 inst_cellmath__24_0_I1108 (.CO(N2441), .S(N2440), .A(N2397), .B(N2430), .CI(N2432));
ADDFHXL inst_cellmath__24_0_I1109 (.CO(N2443), .S(N2442), .A(N2399), .B(N2434), .CI(N2401));
ADDFHXL inst_cellmath__24_0_I1110 (.CO(N2445), .S(N2444), .A(N2438), .B(N2436), .CI(N2403));
ADDFX1 inst_cellmath__24_0_I1111 (.CO(N2447), .S(N2446), .A(N2405), .B(N2440), .CI(N2442));
ADDFHXL inst_cellmath__24_0_I1112 (.CO(N2449), .S(N2448), .A(N2444), .B(N2407), .CI(N2409));
ADDFHXL inst_cellmath__24_0_I1113 (.CO(N2451), .S(N2450), .A(N2411), .B(N2446), .CI(N2448));
ADDFX1 inst_cellmath__24_0_I1114 (.CO(N2453), .S(N2452), .A(N722), .B(N1744), .CI(N779));
ADDFX1 inst_cellmath__24_0_I1115 (.CO(N2455), .S(N2454), .A(N893), .B(N836), .CI(N950));
ADDFX1 inst_cellmath__24_0_I1116 (.CO(N2457), .S(N2456), .A(N1064), .B(N1007), .CI(N1121));
ADDFX1 inst_cellmath__24_0_I1117 (.CO(N2459), .S(N2458), .A(N1235), .B(N1178), .CI(N1292));
ADDFX1 inst_cellmath__24_0_I1118 (.CO(N2461), .S(N2460), .A(N1406), .B(N1349), .CI(N1463));
ADDFX1 inst_cellmath__24_0_I1119 (.CO(N2463), .S(N2462), .A(N1577), .B(N1520), .CI(N1634));
ADDFX1 inst_cellmath__24_0_I1120 (.CO(N2465), .S(N2464), .A(N2415), .B(N1691), .CI(N2417));
ADDFX1 inst_cellmath__24_0_I1121 (.CO(N2467), .S(N2466), .A(N2421), .B(N2419), .CI(N2423));
ADDFX1 inst_cellmath__24_0_I1122 (.CO(N2469), .S(N2468), .A(N2452), .B(N2425), .CI(N2454));
ADDFX1 inst_cellmath__24_0_I1123 (.CO(N2471), .S(N2470), .A(N2458), .B(N2456), .CI(N2460));
ADDFXL inst_cellmath__24_0_I1124 (.CO(N2473), .S(N2472), .A(N2427), .B(N2462), .CI(N2429));
ADDFX1 inst_cellmath__24_0_I1125 (.CO(N2475), .S(N2474), .A(N2464), .B(N2431), .CI(N2466));
ADDFX1 inst_cellmath__24_0_I1126 (.CO(N2477), .S(N2476), .A(N2435), .B(N2433), .CI(N2468));
ADDFXL inst_cellmath__24_0_I1127 (.CO(N2479), .S(N2478), .A(N2437), .B(N2470), .CI(N2472));
ADDFHXL inst_cellmath__24_0_I1128 (.CO(N2481), .S(N2480), .A(N2441), .B(N2439), .CI(N2474));
ADDFX1 inst_cellmath__24_0_I1129 (.CO(N2483), .S(N2482), .A(N2443), .B(N2476), .CI(N2478));
ADDFHXL inst_cellmath__24_0_I1130 (.CO(N2485), .S(N2484), .A(N2480), .B(N2445), .CI(N2447));
ADDFHXL inst_cellmath__24_0_I1131 (.CO(N2487), .S(N2486), .A(N2449), .B(N2482), .CI(N2484));
ADDFX1 inst_cellmath__24_0_I1132 (.CO(N2489), .S(N2488), .A(N781), .B(N1746), .CI(N838));
ADDFX1 inst_cellmath__24_0_I1133 (.CO(N2491), .S(N2490), .A(N952), .B(N895), .CI(N1009));
ADDFX1 inst_cellmath__24_0_I1134 (.CO(N2493), .S(N2492), .A(N1123), .B(N1066), .CI(N1180));
ADDFX1 inst_cellmath__24_0_I1135 (.CO(N2495), .S(N2494), .A(N1294), .B(N1237), .CI(N1351));
ADDFX1 inst_cellmath__24_0_I1136 (.CO(N2497), .S(N2496), .A(N1465), .B(N1408), .CI(N1522));
ADDFX1 inst_cellmath__24_0_I1137 (.CO(N2499), .S(N2498), .A(N1636), .B(N1579), .CI(N1693));
ADDFX1 inst_cellmath__24_0_I1138 (.CO(N2501), .S(N2500), .A(N2455), .B(N2453), .CI(N2457));
ADDFX1 inst_cellmath__24_0_I1139 (.CO(N2503), .S(N2502), .A(N2461), .B(N2459), .CI(N2463));
ADDFX1 inst_cellmath__24_0_I1140 (.CO(N2505), .S(N2504), .A(N2490), .B(N2488), .CI(N2492));
ADDFXL inst_cellmath__24_0_I1141 (.CO(N2507), .S(N2506), .A(N2496), .B(N2494), .CI(N2498));
ADDFX1 inst_cellmath__24_0_I1142 (.CO(N2509), .S(N2508), .A(N2467), .B(N2465), .CI(N2469));
ADDFX1 inst_cellmath__24_0_I1143 (.CO(N2511), .S(N2510), .A(N2500), .B(N2471), .CI(N2502));
ADDFX1 inst_cellmath__24_0_I1144 (.CO(N2513), .S(N2512), .A(N2506), .B(N2473), .CI(N2504));
ADDFHXL inst_cellmath__24_0_I1145 (.CO(N2515), .S(N2514), .A(N2477), .B(N2475), .CI(N2508));
ADDFXL inst_cellmath__24_0_I1146 (.CO(N2517), .S(N2516), .A(N2479), .B(N2510), .CI(N2512));
ADDFHXL inst_cellmath__24_0_I1147 (.CO(N2519), .S(N2518), .A(N2514), .B(N2481), .CI(N2483));
ADDFHXL inst_cellmath__24_0_I1148 (.CO(N2521), .S(N2520), .A(N2485), .B(N2516), .CI(N2518));
ADDFX1 inst_cellmath__24_0_I1149 (.CO(N2523), .S(N2522), .A(N840), .B(N1748), .CI(N897));
ADDFX1 inst_cellmath__24_0_I1150 (.CO(N2525), .S(N2524), .A(N1011), .B(N954), .CI(N1068));
ADDFX1 inst_cellmath__24_0_I1151 (.CO(N2527), .S(N2526), .A(N1182), .B(N1125), .CI(N1239));
ADDFX1 inst_cellmath__24_0_I1152 (.CO(N2529), .S(N2528), .A(N1353), .B(N1296), .CI(N1410));
ADDFX1 inst_cellmath__24_0_I1153 (.CO(N2531), .S(N2530), .A(N1524), .B(N1467), .CI(N1581));
ADDFX1 inst_cellmath__24_0_I1154 (.CO(N2533), .S(N2532), .A(N1695), .B(N1638), .CI(N2489));
ADDFX1 inst_cellmath__24_0_I1155 (.CO(N2535), .S(N2534), .A(N2493), .B(N2491), .CI(N2495));
ADDFX1 inst_cellmath__24_0_I1156 (.CO(N2537), .S(N2536), .A(N2499), .B(N2497), .CI(N2522));
ADDFX1 inst_cellmath__24_0_I1157 (.CO(N2539), .S(N2538), .A(N2526), .B(N2524), .CI(N2528));
ADDFX1 inst_cellmath__24_0_I1158 (.CO(N2541), .S(N2540), .A(N2501), .B(N2530), .CI(N2503));
ADDFX1 inst_cellmath__24_0_I1159 (.CO(N2543), .S(N2542), .A(N2505), .B(N2532), .CI(N2534));
ADDFXL inst_cellmath__24_0_I1160 (.CO(N2545), .S(N2544), .A(N2536), .B(N2507), .CI(N2538));
ADDFX1 inst_cellmath__24_0_I1161 (.CO(N2547), .S(N2546), .A(N2511), .B(N2509), .CI(N2540));
ADDFX1 inst_cellmath__24_0_I1162 (.CO(N2549), .S(N2548), .A(N2513), .B(N2542), .CI(N2544));
ADDFXL inst_cellmath__24_0_I1163 (.CO(N2551), .S(N2550), .A(N2546), .B(N2515), .CI(N2517));
ADDFHXL inst_cellmath__24_0_I1164 (.CO(N2553), .S(N2552), .A(N2519), .B(N2548), .CI(N2550));
ADDFX1 inst_cellmath__24_0_I1165 (.CO(N2555), .S(N2554), .A(N899), .B(N1750), .CI(N956));
ADDFX1 inst_cellmath__24_0_I1166 (.CO(N2557), .S(N2556), .A(N1070), .B(N1013), .CI(N1127));
ADDFX1 inst_cellmath__24_0_I1167 (.CO(N2559), .S(N2558), .A(N1241), .B(N1184), .CI(N1298));
ADDFX1 inst_cellmath__24_0_I1168 (.CO(N2561), .S(N2560), .A(N1412), .B(N1355), .CI(N1469));
ADDFX1 inst_cellmath__24_0_I1169 (.CO(N2563), .S(N2562), .A(N1583), .B(N1526), .CI(N1640));
ADDFX1 inst_cellmath__24_0_I1170 (.CO(N2565), .S(N2564), .A(N2523), .B(N1697), .CI(N2525));
ADDFX1 inst_cellmath__24_0_I1171 (.CO(N2567), .S(N2566), .A(N2529), .B(N2527), .CI(N2531));
ADDFXL inst_cellmath__24_0_I1172 (.CO(N2569), .S(N2568), .A(N2556), .B(N2554), .CI(N2558));
ADDFX1 inst_cellmath__24_0_I1173 (.CO(N2571), .S(N2570), .A(N2562), .B(N2560), .CI(N2533));
ADDFX1 inst_cellmath__24_0_I1174 (.CO(N2573), .S(N2572), .A(N2537), .B(N2535), .CI(N2564));
ADDFXL inst_cellmath__24_0_I1175 (.CO(N2575), .S(N2574), .A(N2566), .B(N2539), .CI(N2568));
ADDFX1 inst_cellmath__24_0_I1176 (.CO(N2577), .S(N2576), .A(N2570), .B(N2541), .CI(N2543));
ADDFX1 inst_cellmath__24_0_I1177 (.CO(N2579), .S(N2578), .A(N2545), .B(N2572), .CI(N2574));
ADDFXL inst_cellmath__24_0_I1178 (.CO(N2581), .S(N2580), .A(N2576), .B(N2547), .CI(N2549));
ADDFX1 inst_cellmath__24_0_I1179 (.CO(N2583), .S(N2582), .A(N2551), .B(N2578), .CI(N2580));
ADDFX1 inst_cellmath__24_0_I1180 (.CO(N2585), .S(N2584), .A(N958), .B(N1752), .CI(N1015));
ADDFX1 inst_cellmath__24_0_I1181 (.CO(N2587), .S(N2586), .A(N1129), .B(N1072), .CI(N1186));
ADDFX1 inst_cellmath__24_0_I1182 (.CO(N2589), .S(N2588), .A(N1300), .B(N1243), .CI(N1357));
ADDFX1 inst_cellmath__24_0_I1183 (.CO(N2591), .S(N2590), .A(N1471), .B(N1414), .CI(N1528));
ADDFX1 inst_cellmath__24_0_I1184 (.CO(N2593), .S(N2592), .A(N1642), .B(N1585), .CI(N1699));
ADDFX1 inst_cellmath__24_0_I1185 (.CO(N2595), .S(N2594), .A(N2557), .B(N2555), .CI(N2559));
ADDFX1 inst_cellmath__24_0_I1186 (.CO(N2597), .S(N2596), .A(N2563), .B(N2561), .CI(N2584));
ADDFX1 inst_cellmath__24_0_I1187 (.CO(N2599), .S(N2598), .A(N2588), .B(N2586), .CI(N2590));
ADDFX1 inst_cellmath__24_0_I1188 (.CO(N2601), .S(N2600), .A(N2565), .B(N2592), .CI(N2567));
ADDFX1 inst_cellmath__24_0_I1189 (.CO(N2603), .S(N2602), .A(N2594), .B(N2569), .CI(N2571));
ADDFX1 inst_cellmath__24_0_I1190 (.CO(N2605), .S(N2604), .A(N2598), .B(N2596), .CI(N2573));
ADDFX1 inst_cellmath__24_0_I1191 (.CO(N2607), .S(N2606), .A(N2575), .B(N2600), .CI(N2602));
ADDFXL inst_cellmath__24_0_I1192 (.CO(N2609), .S(N2608), .A(N2604), .B(N2577), .CI(N2579));
ADDFX1 inst_cellmath__24_0_I1193 (.CO(N2611), .S(N2610), .A(N2581), .B(N2606), .CI(N2608));
ADDFX1 inst_cellmath__24_0_I1194 (.CO(N2613), .S(N2612), .A(N1017), .B(N1754), .CI(N1074));
ADDFX1 inst_cellmath__24_0_I1195 (.CO(N2615), .S(N2614), .A(N1188), .B(N1131), .CI(N1245));
ADDFX1 inst_cellmath__24_0_I1196 (.CO(N2617), .S(N2616), .A(N1359), .B(N1302), .CI(N1416));
ADDFX1 inst_cellmath__24_0_I1197 (.CO(N2619), .S(N2618), .A(N1530), .B(N1473), .CI(N1587));
ADDFX1 inst_cellmath__24_0_I1198 (.CO(N2621), .S(N2620), .A(N1701), .B(N1644), .CI(N2585));
ADDFX1 inst_cellmath__24_0_I1199 (.CO(N2623), .S(N2622), .A(N2589), .B(N2587), .CI(N2591));
ADDFX1 inst_cellmath__24_0_I1200 (.CO(N2625), .S(N2624), .A(N2612), .B(N2593), .CI(N2614));
ADDFX1 inst_cellmath__24_0_I1201 (.CO(N2627), .S(N2626), .A(N2618), .B(N2616), .CI(N2595));
ADDFX1 inst_cellmath__24_0_I1202 (.CO(N2629), .S(N2628), .A(N2620), .B(N2597), .CI(N2599));
ADDFX1 inst_cellmath__24_0_I1203 (.CO(N2631), .S(N2630), .A(N2624), .B(N2622), .CI(N2601));
ADDFX1 inst_cellmath__24_0_I1204 (.CO(N2633), .S(N2632), .A(N2603), .B(N2626), .CI(N2628));
ADDFX1 inst_cellmath__24_0_I1205 (.CO(N2635), .S(N2634), .A(N2630), .B(N2605), .CI(N2607));
ADDFHXL inst_cellmath__24_0_I1206 (.CO(N2637), .S(N2636), .A(N2609), .B(N2632), .CI(N2634));
ADDFX1 inst_cellmath__24_0_I1207 (.CO(N2639), .S(N2638), .A(N1076), .B(N1756), .CI(N1133));
ADDFX1 inst_cellmath__24_0_I1208 (.CO(N2641), .S(N2640), .A(N1247), .B(N1190), .CI(N1304));
ADDFX1 inst_cellmath__24_0_I1209 (.CO(N2643), .S(N2642), .A(N1418), .B(N1361), .CI(N1475));
ADDFX1 inst_cellmath__24_0_I1210 (.CO(N2645), .S(N2644), .A(N1589), .B(N1532), .CI(N1646));
ADDFX1 inst_cellmath__24_0_I1211 (.CO(N2647), .S(N2646), .A(N2613), .B(N1703), .CI(N2615));
ADDFX1 inst_cellmath__24_0_I1212 (.CO(N2649), .S(N2648), .A(N2619), .B(N2617), .CI(N2638));
ADDFX1 inst_cellmath__24_0_I1213 (.CO(N2651), .S(N2650), .A(N2642), .B(N2640), .CI(N2644));
ADDFX1 inst_cellmath__24_0_I1214 (.CO(N2653), .S(N2652), .A(N2623), .B(N2621), .CI(N2625));
ADDFX1 inst_cellmath__24_0_I1215 (.CO(N2655), .S(N2654), .A(N2648), .B(N2646), .CI(N2627));
ADDFX1 inst_cellmath__24_0_I1216 (.CO(N2657), .S(N2656), .A(N2629), .B(N2650), .CI(N2652));
ADDFX1 inst_cellmath__24_0_I1217 (.CO(N2659), .S(N2658), .A(N2654), .B(N2631), .CI(N2633));
ADDFX1 inst_cellmath__24_0_I1218 (.CO(N2661), .S(N2660), .A(N2635), .B(N2656), .CI(N2658));
ADDFX1 inst_cellmath__24_0_I1219 (.CO(N2663), .S(N2662), .A(N1135), .B(N1758), .CI(N1192));
ADDFX1 inst_cellmath__24_0_I1220 (.CO(N2665), .S(N2664), .A(N1306), .B(N1249), .CI(N1363));
ADDFX1 inst_cellmath__24_0_I1221 (.CO(N2667), .S(N2666), .A(N1477), .B(N1420), .CI(N1534));
ADDFX1 inst_cellmath__24_0_I1222 (.CO(N2669), .S(N2668), .A(N1648), .B(N1591), .CI(N1705));
ADDFX1 inst_cellmath__24_0_I1223 (.CO(N2671), .S(N2670), .A(N2641), .B(N2639), .CI(N2643));
ADDFX1 inst_cellmath__24_0_I1224 (.CO(N2673), .S(N2672), .A(N2662), .B(N2645), .CI(N2664));
ADDFX1 inst_cellmath__24_0_I1225 (.CO(N2675), .S(N2674), .A(N2668), .B(N2666), .CI(N2647));
ADDFX1 inst_cellmath__24_0_I1226 (.CO(N2677), .S(N2676), .A(N2651), .B(N2649), .CI(N2670));
ADDFX1 inst_cellmath__24_0_I1227 (.CO(N2679), .S(N2678), .A(N2674), .B(N2672), .CI(N2653));
ADDFX1 inst_cellmath__24_0_I1228 (.CO(N2681), .S(N2680), .A(N2676), .B(N2655), .CI(N2657));
ADDFX1 inst_cellmath__24_0_I1229 (.CO(N2683), .S(N2682), .A(N2659), .B(N2678), .CI(N2680));
ADDFX1 inst_cellmath__24_0_I1230 (.CO(N2685), .S(N2684), .A(N1194), .B(N1760), .CI(N1251));
ADDFX1 inst_cellmath__24_0_I1231 (.CO(N2687), .S(N2686), .A(N1365), .B(N1308), .CI(N1422));
ADDFX1 inst_cellmath__24_0_I1232 (.CO(N2689), .S(N2688), .A(N1536), .B(N1479), .CI(N1593));
ADDFX1 inst_cellmath__24_0_I1233 (.CO(N2691), .S(N2690), .A(N1707), .B(N1650), .CI(N2663));
ADDFX1 inst_cellmath__24_0_I1234 (.CO(N2693), .S(N2692), .A(N2667), .B(N2665), .CI(N2669));
ADDFX1 inst_cellmath__24_0_I1235 (.CO(N2695), .S(N2694), .A(N2686), .B(N2684), .CI(N2688));
ADDFX1 inst_cellmath__24_0_I1236 (.CO(N2697), .S(N2696), .A(N2690), .B(N2671), .CI(N2673));
ADDFX1 inst_cellmath__24_0_I1237 (.CO(N2699), .S(N2698), .A(N2675), .B(N2692), .CI(N2694));
ADDFX1 inst_cellmath__24_0_I1238 (.CO(N2701), .S(N2700), .A(N2696), .B(N2677), .CI(N2679));
ADDFX1 inst_cellmath__24_0_I1239 (.CO(N2703), .S(N2702), .A(N2681), .B(N2698), .CI(N2700));
ADDFX1 inst_cellmath__24_0_I1240 (.CO(N2705), .S(N2704), .A(N1253), .B(N1762), .CI(N1310));
ADDFX1 inst_cellmath__24_0_I1241 (.CO(N2707), .S(N2706), .A(N1424), .B(N1367), .CI(N1481));
ADDFX1 inst_cellmath__24_0_I1242 (.CO(N2709), .S(N2708), .A(N1595), .B(N1538), .CI(N1652));
ADDFX1 inst_cellmath__24_0_I1243 (.CO(N2711), .S(N2710), .A(N2685), .B(N1709), .CI(N2687));
ADDFX1 inst_cellmath__24_0_I1244 (.CO(N2713), .S(N2712), .A(N2704), .B(N2689), .CI(N2706));
ADDFX1 inst_cellmath__24_0_I1245 (.CO(N2715), .S(N2714), .A(N2691), .B(N2708), .CI(N2693));
ADDFX1 inst_cellmath__24_0_I1246 (.CO(N2717), .S(N2716), .A(N2695), .B(N2710), .CI(N2712));
ADDFX1 inst_cellmath__24_0_I1247 (.CO(N2719), .S(N2718), .A(N2714), .B(N2697), .CI(N2699));
ADDFX1 inst_cellmath__24_0_I1248 (.CO(N2721), .S(N2720), .A(N2701), .B(N2716), .CI(N2718));
ADDFX1 inst_cellmath__24_0_I1249 (.CO(N2723), .S(N2722), .A(N1312), .B(N1764), .CI(N1369));
ADDFX1 inst_cellmath__24_0_I1250 (.CO(N2725), .S(N2724), .A(N1483), .B(N1426), .CI(N1540));
ADDFX1 inst_cellmath__24_0_I1251 (.CO(N2727), .S(N2726), .A(N1654), .B(N1597), .CI(N1711));
ADDFX1 inst_cellmath__24_0_I1252 (.CO(N2729), .S(N2728), .A(N2707), .B(N2705), .CI(N2709));
ADDFX1 inst_cellmath__24_0_I1253 (.CO(N2731), .S(N2730), .A(N2724), .B(N2722), .CI(N2726));
ADDFX1 inst_cellmath__24_0_I1254 (.CO(N2733), .S(N2732), .A(N2713), .B(N2711), .CI(N2728));
ADDFX1 inst_cellmath__24_0_I1255 (.CO(N2735), .S(N2734), .A(N2730), .B(N2715), .CI(N2717));
ADDFX1 inst_cellmath__24_0_I1256 (.CO(N2737), .S(N2736), .A(N2719), .B(N2732), .CI(N2734));
ADDFX1 inst_cellmath__24_0_I1257 (.CO(N2739), .S(N2738), .A(N1371), .B(N1766), .CI(N1428));
ADDFX1 inst_cellmath__24_0_I1258 (.CO(N2741), .S(N2740), .A(N1542), .B(N1485), .CI(N1599));
ADDFX1 inst_cellmath__24_0_I1259 (.CO(N2743), .S(N2742), .A(N1713), .B(N1656), .CI(N2723));
ADDFX1 inst_cellmath__24_0_I1260 (.CO(N2745), .S(N2744), .A(N2727), .B(N2725), .CI(N2738));
ADDFX1 inst_cellmath__24_0_I1261 (.CO(N2747), .S(N2746), .A(N2729), .B(N2740), .CI(N2742));
ADDFX1 inst_cellmath__24_0_I1262 (.CO(N2749), .S(N2748), .A(N2744), .B(N2731), .CI(N2733));
ADDFX1 inst_cellmath__24_0_I1263 (.CO(N2751), .S(N2750), .A(N2735), .B(N2746), .CI(N2748));
ADDFX1 inst_cellmath__24_0_I1264 (.CO(N2753), .S(N2752), .A(N1430), .B(N1768), .CI(N1487));
ADDFX1 inst_cellmath__24_0_I1265 (.CO(N2755), .S(N2754), .A(N1601), .B(N1544), .CI(N1658));
ADDFX1 inst_cellmath__24_0_I1266 (.CO(N2757), .S(N2756), .A(N2739), .B(N1715), .CI(N2741));
ADDFX1 inst_cellmath__24_0_I1267 (.CO(N2759), .S(N2758), .A(N2754), .B(N2752), .CI(N2743));
ADDFX1 inst_cellmath__24_0_I1268 (.CO(N2761), .S(N2760), .A(N2756), .B(N2745), .CI(N2747));
ADDFX1 inst_cellmath__24_0_I1269 (.CO(N2763), .S(N2762), .A(N2749), .B(N2758), .CI(N2760));
ADDFX1 inst_cellmath__24_0_I1270 (.CO(N2765), .S(N2764), .A(N1489), .B(N1770), .CI(N1546));
ADDFX1 inst_cellmath__24_0_I1271 (.CO(N2767), .S(N2766), .A(N1660), .B(N1603), .CI(N1717));
ADDFX1 inst_cellmath__24_0_I1272 (.CO(N2769), .S(N2768), .A(N2755), .B(N2753), .CI(N2764));
ADDFX1 inst_cellmath__24_0_I1273 (.CO(N2771), .S(N2770), .A(N2757), .B(N2766), .CI(N2759));
ADDFX1 inst_cellmath__24_0_I1274 (.CO(N2773), .S(N2772), .A(N2761), .B(N2768), .CI(N2770));
ADDFX1 inst_cellmath__24_0_I1275 (.CO(N2775), .S(N2774), .A(N1548), .B(N1772), .CI(N1605));
ADDFX1 inst_cellmath__24_0_I1276 (.CO(N2777), .S(N2776), .A(N1719), .B(N1662), .CI(N2765));
ADDFX1 inst_cellmath__24_0_I1277 (.CO(N2779), .S(N2778), .A(N2774), .B(N2767), .CI(N2769));
ADDFX1 inst_cellmath__24_0_I1278 (.CO(N2781), .S(N2780), .A(N2771), .B(N2776), .CI(N2778));
ADDFX1 inst_cellmath__24_0_I1279 (.CO(N2783), .S(N2782), .A(N1607), .B(N1774), .CI(N1664));
ADDFX1 inst_cellmath__24_0_I1280 (.CO(N2785), .S(N2784), .A(N2775), .B(N1721), .CI(N2782));
ADDFX1 inst_cellmath__24_0_I1281 (.CO(N2787), .S(N2786), .A(N2784), .B(N2777), .CI(N2779));
ADDFX1 inst_cellmath__24_0_I1282 (.CO(N2789), .S(N2788), .A(N1666), .B(N1776), .CI(N1723));
ADDFX1 inst_cellmath__24_0_I1283 (.CO(N2791), .S(N2790), .A(N2788), .B(N2783), .CI(N2785));
ADDFX1 inst_cellmath__24_0_I1284 (.CO(N3110), .S(N2792), .A(N1725), .B(N1778), .CI(N2789));
NAND2XL inst_cellmath__24_0_I1285 (.Y(N2794), .A(N383), .B(N440));
NOR2XL inst_cellmath__24_0_I1286 (.Y(N2795), .A(N499), .B(N1782));
NAND2XL inst_cellmath__24_0_I1287 (.Y(N2796), .A(N499), .B(N1782));
NOR2XL inst_cellmath__24_0_I1288 (.Y(N2797), .A(N1784), .B(N1786));
NAND2XL inst_cellmath__24_0_I1289 (.Y(N2798), .A(N1784), .B(N1786));
NOR2XL inst_cellmath__24_0_I1290 (.Y(N2799), .A(N1787), .B(N1792));
NAND2XL inst_cellmath__24_0_I1291 (.Y(N2800), .A(N1787), .B(N1792));
NOR2XL inst_cellmath__24_0_I1292 (.Y(N2801), .A(N1798), .B(N1800));
NAND2XL inst_cellmath__24_0_I1293 (.Y(N2802), .A(N1798), .B(N1800));
NOR2XL inst_cellmath__24_0_I1294 (.Y(N2803), .A(N1801), .B(N1810));
NAND2XL inst_cellmath__24_0_I1295 (.Y(N2804), .A(N1801), .B(N1810));
NOR2XL inst_cellmath__24_0_I1296 (.Y(N2805), .A(N1811), .B(N1822));
NAND2XL inst_cellmath__24_0_I1297 (.Y(N2806), .A(N1811), .B(N1822));
NOR2X1 inst_cellmath__24_0_I1298 (.Y(N2807), .A(N1823), .B(N1836));
NAND2XL inst_cellmath__24_0_I1299 (.Y(N2808), .A(N1823), .B(N1836));
NOR2XL inst_cellmath__24_0_I1300 (.Y(N2809), .A(N1837), .B(N1852));
NAND2X1 inst_cellmath__24_0_I1301 (.Y(N2810), .A(N1837), .B(N1852));
NOR2X2 inst_cellmath__24_0_I1302 (.Y(N2811), .A(N1853), .B(N1870));
NAND2X1 inst_cellmath__24_0_I1303 (.Y(N2812), .A(N1853), .B(N1870));
NOR2XL inst_cellmath__24_0_I1304 (.Y(N2813), .A(N1871), .B(N1890));
NAND2X2 inst_cellmath__24_0_I1305 (.Y(N2814), .A(N1871), .B(N1890));
NOR2XL inst_cellmath__24_0_I1306 (.Y(N2815), .A(N1891), .B(N1912));
NAND2XL inst_cellmath__24_0_I1307 (.Y(N2816), .A(N1891), .B(N1912));
NOR2X1 inst_cellmath__24_0_I1308 (.Y(N2817), .A(N1913), .B(N1936));
NAND2XL inst_cellmath__24_0_I1309 (.Y(N2818), .A(N1913), .B(N1936));
NOR2XL inst_cellmath__24_0_I1310 (.Y(N2819), .A(N1937), .B(N1962));
NAND2X2 inst_cellmath__24_0_I1311 (.Y(N2820), .A(N1937), .B(N1962));
AOI21XL inst_cellmath__24_0_I1314 (.Y(N2823), .A0(N2796), .A1(N2794), .B0(N2795));
INVXL inst_cellmath__24_0_I2422 (.Y(N4152), .A(N2797));
INVXL inst_cellmath__24_0_I2423 (.Y(N4153), .A(N2798));
OAI21XL inst_cellmath__24_0_I1322 (.Y(N2831), .A0(N4153), .A1(N2823), .B0(N4152));
AOI21XL inst_cellmath__24_0_I1330 (.Y(N2839), .A0(N2800), .A1(N2831), .B0(N2799));
INVXL inst_cellmath__24_0_I2429 (.Y(N4159), .A(N2801));
INVXL inst_cellmath__24_0_I2430 (.Y(N4160), .A(N2802));
OAI21XL inst_cellmath__24_0_I1342 (.Y(N2851), .A0(N4160), .A1(N2839), .B0(N4159));
AOI21X1 inst_cellmath__24_0_I1354 (.Y(N2863), .A0(N2804), .A1(N2851), .B0(N2803));
INVXL inst_cellmath__24_0_I2440 (.Y(N4170), .A(N2805));
INVXL inst_cellmath__24_0_I2441 (.Y(N4171), .A(N2806));
OAI21X1 inst_cellmath__24_0_I1370 (.Y(N2879), .A0(N4171), .A1(N2863), .B0(N4170));
AO21XL inst_cellmath__24_0_I2812 (.Y(N4182), .A0(N2810), .A1(N2807), .B0(N2809));
CLKAND2X2 inst_cellmath__24_0_I2683 (.Y(N4183), .A(N2810), .B(N2808));
AOI21XL inst_cellmath__24_0_I1394 (.Y(N2903), .A0(N2808), .A1(N2879), .B0(N2807));
AOI21X2 inst_cellmath__24_0_I1396 (.Y(N2905), .A0(N4183), .A1(N2879), .B0(N4182));
AOI21X2 inst_cellmath__24_0_I1400 (.Y(N2909), .A0(N2814), .A1(N2811), .B0(N2813));
NAND2X2 inst_cellmath__24_0_I1401 (.Y(N2910), .A(N2814), .B(N2812));
OAI21X2 inst_cellmath__24_0_I1422 (.Y(N2931), .A0(N2910), .A1(N2905), .B0(N2909));
NOR2BX1 andori2bb1_A_I6135 (.Y(N4346), .AN(N2812), .B(N2905));
NOR2XL andori2bb1_A_I2852 (.Y(N4213), .A(N4346), .B(N2811));
AOI21X2 inst_cellmath__24_0_I1446 (.Y(N2955), .A0(N2816), .A1(N2931), .B0(N2815));
INVXL inst_cellmath__24_0_I2487 (.Y(N4217), .A(N2817));
INVXL inst_cellmath__24_0_I2488 (.Y(N4218), .A(N2818));
AOI21X2 inst_cellmath__24_0_I1450 (.Y(N2959), .A0(N2820), .A1(N2817), .B0(N2819));
NAND2X1 inst_cellmath__24_0_I1451 (.Y(N2960), .A(N2820), .B(N2818));
OAI21XL inst_cellmath__24_0_I1476 (.Y(N2985), .A0(N4218), .A1(N2955), .B0(N4217));
OAI21X2 inst_cellmath__24_0_I1478 (.Y(N3046), .A0(N2960), .A1(N2955), .B0(N2959));
NAND2BXL inst_cellmath__24_0_I1485 (.Y(N2994), .AN(N2795), .B(N2796));
NAND2BXL inst_cellmath__24_0_I1488 (.Y(N2997), .AN(N2797), .B(N2798));
NAND2BXL inst_cellmath__24_0_I1491 (.Y(N3000), .AN(N2799), .B(N2800));
NAND2BXL inst_cellmath__24_0_I1494 (.Y(N3003), .AN(N2801), .B(N2802));
NAND2BXL inst_cellmath__24_0_I1497 (.Y(N3006), .AN(N2803), .B(N2804));
NAND2BXL inst_cellmath__24_0_I1500 (.Y(N3009), .AN(N2805), .B(N2806));
NAND2BXL inst_cellmath__24_0_I1503 (.Y(N3012), .AN(N2807), .B(N2808));
NAND2BXL inst_cellmath__24_0_I1506 (.Y(N3015), .AN(N2809), .B(N2810));
NAND2BXL inst_cellmath__24_0_I1509 (.Y(N3018), .AN(N2811), .B(N2812));
NAND2BXL inst_cellmath__24_0_I1512 (.Y(N3021), .AN(N2813), .B(N2814));
NAND2BXL inst_cellmath__24_0_I1515 (.Y(N3024), .AN(N2815), .B(N2816));
NAND2BXL inst_cellmath__24_0_I1518 (.Y(N3027), .AN(N2817), .B(N2818));
NAND2BXL inst_cellmath__24_0_I1521 (.Y(N3030), .AN(N2819), .B(N2820));
XOR2XL inst_cellmath__24_0_I1522 (.Y(inst_cellmath__24_0_out0[1]), .A(N383), .B(N440));
XOR2XL inst_cellmath__24_0_I2687 (.Y(inst_cellmath__24_0_out0[2]), .A(N2794), .B(N2994));
XNOR2X1 inst_cellmath__24_0_I1524 (.Y(inst_cellmath__24_0_out0[3]), .A(N2823), .B(N2997));
XOR2XL inst_cellmath__24_0_I2688 (.Y(inst_cellmath__24_0_out0[4]), .A(N2831), .B(N3000));
XNOR2X1 inst_cellmath__24_0_I1526 (.Y(inst_cellmath__24_0_out0[5]), .A(N2839), .B(N3003));
XOR2XL inst_cellmath__24_0_I2689 (.Y(inst_cellmath__24_0_out0[6]), .A(N2851), .B(N3006));
XNOR2X1 inst_cellmath__24_0_I1528 (.Y(inst_cellmath__24_0_out0[7]), .A(N2863), .B(N3009));
XOR2XL inst_cellmath__24_0_I2690 (.Y(inst_cellmath__24_0_out0[8]), .A(N2879), .B(N3012));
XNOR2X1 inst_cellmath__24_0_I1530 (.Y(inst_cellmath__24_0_out0[9]), .A(N2903), .B(N3015));
XNOR2X1 inst_cellmath__24_0_I1531 (.Y(inst_cellmath__24_0_out0[10]), .A(N2905), .B(N3018));
XNOR2X1 inst_cellmath__24_0_I1532 (.Y(inst_cellmath__24_0_out0[11]), .A(N4213), .B(N3021));
XOR2XL inst_cellmath__24_0_I2691 (.Y(inst_cellmath__24_0_out0[12]), .A(N2931), .B(N3024));
XNOR2X1 inst_cellmath__24_0_I1534 (.Y(inst_cellmath__24_0_out0[13]), .A(N2955), .B(N3027));
XOR2XL inst_cellmath__24_0_I1535 (.Y(inst_cellmath__24_0_out0[14]), .A(N2985), .B(N3030));
NOR2XL inst_cellmath__24_0_I1538 (.Y(N3048), .A(N1963), .B(N1990));
NAND2XL inst_cellmath__24_0_I1539 (.Y(N3049), .A(N1963), .B(N1990));
NOR2X2 inst_cellmath__24_0_I1540 (.Y(N3050), .A(N1991), .B(N2020));
NAND2X1 inst_cellmath__24_0_I1541 (.Y(N3051), .A(N1991), .B(N2020));
NOR2X1 inst_cellmath__24_0_I1542 (.Y(N3052), .A(N2021), .B(N2052));
NAND2X4 inst_cellmath__24_0_I1543 (.Y(N3053), .A(N2021), .B(N2052));
NOR2X1 inst_cellmath__24_0_I1544 (.Y(N3054), .A(N2053), .B(N2086));
NAND2X2 inst_cellmath__24_0_I1545 (.Y(N3055), .A(N2053), .B(N2086));
NOR2XL inst_cellmath__24_0_I1546 (.Y(N3056), .A(N2087), .B(N2122));
NAND2X4 inst_cellmath__24_0_I1547 (.Y(N3057), .A(N2087), .B(N2122));
NOR2X2 inst_cellmath__24_0_I1548 (.Y(N3058), .A(N2123), .B(N2160));
NAND2X1 inst_cellmath__24_0_I1549 (.Y(N3059), .A(N2123), .B(N2160));
NOR2X1 inst_cellmath__24_0_I1550 (.Y(N3060), .A(N2161), .B(N2200));
NAND2X2 inst_cellmath__24_0_I1551 (.Y(N3061), .A(N2161), .B(N2200));
NOR2X2 inst_cellmath__24_0_I1552 (.Y(N3062), .A(N2201), .B(N2242));
NAND2X2 inst_cellmath__24_0_I1553 (.Y(N3063), .A(N2201), .B(N2242));
NOR2X1 inst_cellmath__24_0_I1554 (.Y(N3064), .A(N2243), .B(N2286));
NAND2X4 inst_cellmath__24_0_I1555 (.Y(N3065), .A(N2243), .B(N2286));
NOR2X2 inst_cellmath__24_0_I1556 (.Y(N3066), .A(N2287), .B(N2330));
NAND2XL inst_cellmath__24_0_I1557 (.Y(N3067), .A(N2287), .B(N2330));
NOR2XL inst_cellmath__24_0_I1558 (.Y(N3068), .A(N2331), .B(N2372));
NAND2X2 inst_cellmath__24_0_I1559 (.Y(N3069), .A(N2331), .B(N2372));
NOR2X2 inst_cellmath__24_0_I1560 (.Y(N3070), .A(N2373), .B(N2412));
NAND2X2 inst_cellmath__24_0_I1561 (.Y(N3071), .A(N2373), .B(N2412));
NOR2XL inst_cellmath__24_0_I1562 (.Y(N3072), .A(N2413), .B(N2450));
NAND2X4 inst_cellmath__24_0_I1563 (.Y(N3073), .A(N2413), .B(N2450));
NOR2X2 inst_cellmath__24_0_I1564 (.Y(N3074), .A(N2451), .B(N2486));
NAND2X2 inst_cellmath__24_0_I1565 (.Y(N3075), .A(N2451), .B(N2486));
NOR2X1 inst_cellmath__24_0_I1566 (.Y(N3076), .A(N2487), .B(N2520));
NAND2X4 inst_cellmath__24_0_I1567 (.Y(N3077), .A(N2487), .B(N2520));
NOR2X1 inst_cellmath__24_0_I1568 (.Y(N3078), .A(N2521), .B(N2552));
NAND2X2 inst_cellmath__24_0_I1569 (.Y(N3079), .A(N2521), .B(N2552));
NOR2XL inst_cellmath__24_0_I1570 (.Y(N3080), .A(N2553), .B(N2582));
NAND2X4 inst_cellmath__24_0_I1571 (.Y(N3081), .A(N2553), .B(N2582));
NOR2X2 inst_cellmath__24_0_I1572 (.Y(N3082), .A(N2583), .B(N2610));
NAND2X1 inst_cellmath__24_0_I1573 (.Y(N3083), .A(N2583), .B(N2610));
NOR2X1 inst_cellmath__24_0_I1574 (.Y(N3084), .A(N2611), .B(N2636));
NAND2X4 inst_cellmath__24_0_I1575 (.Y(N3085), .A(N2611), .B(N2636));
NOR2X1 inst_cellmath__24_0_I1576 (.Y(N3086), .A(N2637), .B(N2660));
NAND2X1 inst_cellmath__24_0_I1577 (.Y(N3087), .A(N2637), .B(N2660));
NOR2XL inst_cellmath__24_0_I1578 (.Y(N3088), .A(N2661), .B(N2682));
NAND2X2 inst_cellmath__24_0_I1579 (.Y(N3089), .A(N2661), .B(N2682));
NOR2XL inst_cellmath__24_0_I1580 (.Y(N3090), .A(N2683), .B(N2702));
NAND2XL inst_cellmath__24_0_I1581 (.Y(N3091), .A(N2683), .B(N2702));
NOR2XL inst_cellmath__24_0_I1582 (.Y(N3092), .A(N2703), .B(N2720));
NAND2XL inst_cellmath__24_0_I1583 (.Y(N3093), .A(N2703), .B(N2720));
NOR2XL inst_cellmath__24_0_I1584 (.Y(N3094), .A(N2721), .B(N2736));
NAND2XL inst_cellmath__24_0_I1585 (.Y(N3095), .A(N2721), .B(N2736));
NOR2XL inst_cellmath__24_0_I1586 (.Y(N3096), .A(N2737), .B(N2750));
NAND2XL inst_cellmath__24_0_I1587 (.Y(N3097), .A(N2737), .B(N2750));
NOR2XL inst_cellmath__24_0_I1588 (.Y(N3098), .A(N2751), .B(N2762));
NAND2XL inst_cellmath__24_0_I1589 (.Y(N3099), .A(N2751), .B(N2762));
NOR2XL inst_cellmath__24_0_I1590 (.Y(N3100), .A(N2763), .B(N2772));
NAND2XL inst_cellmath__24_0_I1591 (.Y(N3101), .A(N2763), .B(N2772));
NOR2XL inst_cellmath__24_0_I1592 (.Y(N3102), .A(N2773), .B(N2780));
NAND2XL inst_cellmath__24_0_I1593 (.Y(N3103), .A(N2773), .B(N2780));
NOR2XL inst_cellmath__24_0_I1594 (.Y(N3104), .A(N2786), .B(N2781));
NAND2XL inst_cellmath__24_0_I1595 (.Y(N3105), .A(N2786), .B(N2781));
NOR2XL inst_cellmath__24_0_I1596 (.Y(N3106), .A(N2790), .B(N2787));
NAND2XL inst_cellmath__24_0_I1597 (.Y(N3107), .A(N2790), .B(N2787));
NOR2XL inst_cellmath__24_0_I1598 (.Y(N3108), .A(N2792), .B(N2791));
NAND2XL inst_cellmath__24_0_I1599 (.Y(N3109), .A(N2792), .B(N2791));
AOI21X2 inst_cellmath__24_0_I1603 (.Y(N3113), .A0(N3049), .A1(N3046), .B0(N3048));
AOI21X4 inst_cellmath__24_0_I1607 (.Y(N3117), .A0(N3053), .A1(N3050), .B0(N3052));
NAND2X2 inst_cellmath__24_0_I1608 (.Y(N3118), .A(N3053), .B(N3051));
INVXL inst_cellmath__24_0_I2494 (.Y(N4224), .A(N3054));
INVXL inst_cellmath__24_0_I2495 (.Y(N4225), .A(N3055));
AOI21X2 inst_cellmath__24_0_I1611 (.Y(N3121), .A0(N3057), .A1(N3054), .B0(N3056));
NAND2X4 inst_cellmath__24_0_I1612 (.Y(N3122), .A(N3057), .B(N3055));
INVXL inst_cellmath__24_0_I2498 (.Y(N4228), .A(N3117));
OAI21XL inst_cellmath__24_0_I1617 (.Y(N3127), .A0(N4225), .A1(N3117), .B0(N4224));
OAI21X2 inst_cellmath__24_0_I1619 (.Y(N3129), .A0(N3122), .A1(N3117), .B0(N3121));
NOR2X2 inst_cellmath__24_0_I1620 (.Y(N3130), .A(N3122), .B(N3118));
AOI21X2 inst_cellmath__24_0_I1623 (.Y(N3133), .A0(N3061), .A1(N3058), .B0(N3060));
AOI21X4 inst_cellmath__24_0_I1627 (.Y(N3137), .A0(N3065), .A1(N3062), .B0(N3064));
NAND2X4 inst_cellmath__24_0_I1628 (.Y(N3138), .A(N3065), .B(N3063));
AOI21X2 inst_cellmath__24_0_I1631 (.Y(N3141), .A0(N3069), .A1(N3066), .B0(N3068));
AOI21X2 inst_cellmath__24_0_I1635 (.Y(N3145), .A0(N3073), .A1(N3070), .B0(N3072));
NAND2X2 inst_cellmath__24_0_I1636 (.Y(N3146), .A(N3073), .B(N3071));
AOI21X4 inst_cellmath__24_0_I1639 (.Y(N3149), .A0(N3077), .A1(N3074), .B0(N3076));
AOI21X2 inst_cellmath__24_0_I1643 (.Y(N3153), .A0(N3081), .A1(N3078), .B0(N3080));
AOI21X4 inst_cellmath__24_0_I1647 (.Y(N3157), .A0(N3085), .A1(N3082), .B0(N3084));
NAND2X2 inst_cellmath__24_0_I1648 (.Y(N3158), .A(N3085), .B(N3083));
INVXL inst_cellmath__24_0_I2514 (.Y(N4244), .A(N3086));
INVXL inst_cellmath__24_0_I2515 (.Y(N4245), .A(N3087));
AOI21X2 inst_cellmath__24_0_I1651 (.Y(N3161), .A0(N3089), .A1(N3086), .B0(N3088));
NAND2X2 inst_cellmath__24_0_I1652 (.Y(N3162), .A(N3089), .B(N3087));
INVXL inst_cellmath__24_0_I2518 (.Y(N4248), .A(N3157));
OAI21XL inst_cellmath__24_0_I1657 (.Y(N3167), .A0(N4245), .A1(N3157), .B0(N4244));
OAI21X4 inst_cellmath__24_0_I1659 (.Y(N3169), .A0(N3162), .A1(N3157), .B0(N3161));
NOR2X2 inst_cellmath__24_0_I1660 (.Y(N3170), .A(N3162), .B(N3158));
AOI21X1 inst_cellmath__24_0_I1663 (.Y(N3173), .A0(N3093), .A1(N3090), .B0(N3092));
NAND2X1 inst_cellmath__24_0_I1664 (.Y(N3174), .A(N3093), .B(N3091));
INVXL inst_cellmath__24_0_I2522 (.Y(N4252), .A(N3094));
INVXL inst_cellmath__24_0_I2523 (.Y(N4253), .A(N3095));
AOI21XL inst_cellmath__24_0_I1667 (.Y(N3177), .A0(N3097), .A1(N3094), .B0(N3096));
NAND2XL inst_cellmath__24_0_I1668 (.Y(N3178), .A(N3097), .B(N3095));
INVXL inst_cellmath__24_0_I2526 (.Y(N4256), .A(N3173));
OAI21XL inst_cellmath__24_0_I1673 (.Y(N3183), .A0(N4253), .A1(N3173), .B0(N4252));
OAI21X1 inst_cellmath__24_0_I1675 (.Y(N3185), .A0(N3178), .A1(N3173), .B0(N3177));
NOR2X2 inst_cellmath__24_0_I1676 (.Y(N3186), .A(N3178), .B(N3174));
AOI21XL inst_cellmath__24_0_I1679 (.Y(N3189), .A0(N3101), .A1(N3098), .B0(N3100));
NAND2XL inst_cellmath__24_0_I1680 (.Y(N3190), .A(N3101), .B(N3099));
INVXL inst_cellmath__24_0_I2530 (.Y(N4260), .A(N3102));
INVXL inst_cellmath__24_0_I2531 (.Y(N4261), .A(N3103));
AOI21XL inst_cellmath__24_0_I1683 (.Y(N3193), .A0(N3105), .A1(N3102), .B0(N3104));
NAND2XL inst_cellmath__24_0_I1684 (.Y(N3194), .A(N3105), .B(N3103));
INVXL inst_cellmath__24_0_I2534 (.Y(N4264), .A(N3189));
OAI21XL inst_cellmath__24_0_I1689 (.Y(N3199), .A0(N4261), .A1(N3189), .B0(N4260));
AOI21XL inst_cellmath__24_0_I1695 (.Y(N3205), .A0(N3109), .A1(N3106), .B0(N3108));
NAND2XL inst_cellmath__24_0_I1696 (.Y(N3206), .A(N3109), .B(N3107));
INVXL inst_cellmath__24_0_I2542 (.Y(N4272), .A(N3205));
NOR2XL inst_cellmath__24_0_I1703 (.Y(N3505), .A(N3110), .B(N3205));
NOR2XL inst_cellmath__24_0_I1704 (.Y(N3215), .A(N3110), .B(N3206));
INVX2 inst_cellmath__24_0_I2544 (.Y(N4274), .A(N3113));
INVX2 inst_cellmath__24_0_I2547 (.Y(N4277), .A(N3133));
CLKAND2X2 inst_cellmath__24_0_I2695 (.Y(N4278), .A(N3061), .B(N3059));
INVX3 inst_cellmath__24_0_I2551 (.Y(N4281), .A(N3137));
INVX3 inst_cellmath__24_0_I2552 (.Y(N4282), .A(N3138));
INVX3 inst_cellmath__24_0_I2555 (.Y(N4285), .A(N3141));
CLKAND2X2 inst_cellmath__24_0_I2638 (.Y(N4286), .A(N3069), .B(N3067));
INVX2 inst_cellmath__24_0_I2559 (.Y(N4289), .A(N3145));
INVX3 inst_cellmath__24_0_I2560 (.Y(N4290), .A(N3146));
INVX3 inst_cellmath__24_0_I2563 (.Y(N4293), .A(N3149));
CLKAND2X3 inst_cellmath__24_0_I2703 (.Y(N4294), .A(N3077), .B(N3075));
INVX2 inst_cellmath__24_0_I2567 (.Y(N4297), .A(N3153));
CLKAND2X6 inst_cellmath__24_0_I2705 (.Y(N4298), .A(N3081), .B(N3079));
INVXL inst_cellmath__24_0_I2569 (.Y(N4299), .A(N4274));
AOI21X4 inst_cellmath__24_0_I1735 (.Y(N3246), .A0(N3130), .A1(N4274), .B0(N3129));
INVXL inst_cellmath__24_0_I2573 (.Y(N4303), .A(N4278));
AOI21X4 inst_cellmath__24_0_I1739 (.Y(N3250), .A0(N4282), .A1(N4277), .B0(N4281));
NAND2X4 inst_cellmath__24_0_I1740 (.Y(N3251), .A(N4282), .B(N4278));
OAI21X4 inst_cellmath__24_0_I1747 (.Y(N3258), .A0(N3251), .A1(N3246), .B0(N3250));
AOI21X4 inst_cellmath__24_0_I1751 (.Y(N3262), .A0(N4290), .A1(N4285), .B0(N4289));
NAND2X4 inst_cellmath__24_0_I1752 (.Y(N3263), .A(N4290), .B(N4286));
INVXL inst_cellmath__24_0_I2584 (.Y(N4314), .A(N4293));
INVXL inst_cellmath__24_0_I2585 (.Y(N4315), .A(N4294));
AOI21X4 inst_cellmath__24_0_I1755 (.Y(N3266), .A0(N4298), .A1(N4293), .B0(N4297));
NAND2X8 inst_cellmath__24_0_I1756 (.Y(N3267), .A(N4298), .B(N4294));
INVXL inst_cellmath__24_0_I2588 (.Y(N4318), .A(N3262));
INVXL inst_cellmath__24_0_I2589 (.Y(N4319), .A(N3263));
OAI21XL inst_cellmath__24_0_I1761 (.Y(N3272), .A0(N4315), .A1(N3262), .B0(N4314));
NOR2XL inst_cellmath__24_0_I1762 (.Y(N3273), .A(N4315), .B(N3263));
OAI21X4 inst_cellmath__24_0_I1763 (.Y(N3274), .A0(N3267), .A1(N3262), .B0(N3266));
NOR2X4 inst_cellmath__24_0_I1764 (.Y(N3275), .A(N3267), .B(N3263));
NOR2XL andori2bb1_A_I2871 (.Y(N4407), .A(N4303), .B(N3246));
NOR2XL andori2bb1_A_I2872 (.Y(N4322), .A(N4407), .B(N4277));
INVXL inst_cellmath__24_0_I2593 (.Y(N4323), .A(N3258));
AOI21XL inst_cellmath__24_0_I2712 (.Y(N3284), .A0(N4286), .A1(N3258), .B0(N4285));
AOI21XL inst_cellmath__24_0_I1775 (.Y(N3286), .A0(N4319), .A1(N3258), .B0(N4318));
AOI21XL inst_cellmath__24_0_I1777 (.Y(N3288), .A0(N3273), .A1(N3258), .B0(N3272));
AOI21X4 inst_cellmath__24_0_I1779 (.Y(N3290), .A0(N3275), .A1(N3258), .B0(N3274));
INVXL buf1_A_I6164 (.Y(N8767), .A(N3290));
INVXL buf1_A_I6165 (.Y(N4325), .A(N8767));
AOI21X4 inst_cellmath__24_0_I1783 (.Y(N3294), .A0(N3186), .A1(N3169), .B0(N3185));
NAND2X1 inst_cellmath__24_0_I1784 (.Y(N3295), .A(N3186), .B(N3170));
OA21X1 inst_cellmath__24_0_I2714 (.Y(N4328), .A0(N3194), .A1(N3189), .B0(N3193));
OR2XL inst_cellmath__24_0_I2715 (.Y(N4329), .A(N3194), .B(N3190));
OAI21X2 inst_cellmath__24_0_I1791 (.Y(N3302), .A0(N4329), .A1(N3294), .B0(N4328));
INVXL inst_cellmath__24_0_I2604 (.Y(N4334), .A(N3169));
INVXL inst_cellmath__24_0_I2605 (.Y(N4335), .A(N3170));
INVX2 inst_cellmath__24_0_I2608 (.Y(N4338), .A(N3302));
OR2XL inst_cellmath__24_0_I2760 (.Y(N4339), .A(N4329), .B(N3295));
OAI21XL inst_cellmath__24_0_I1815 (.Y(N3326), .A0(N4335), .A1(N4325), .B0(N4334));
OAI21XL inst_cellmath__24_0_I2824 (.Y(N3328), .A0(N3295), .A1(N4325), .B0(N3294));
OAI21X4 inst_cellmath__24_0_I1819 (.Y(N3330), .A0(N4339), .A1(N3290), .B0(N4338));
INVXL inst_cellmath__24_0_I2614 (.Y(N4344), .A(N3330));
NAND2BXL inst_cellmath__24_0_I1826 (.Y(N3337), .AN(N3048), .B(N3049));
NAND2BXL inst_cellmath__24_0_I1829 (.Y(N3340), .AN(N3050), .B(N3051));
NAND2BXL inst_cellmath__24_0_I1832 (.Y(N3343), .AN(N3052), .B(N3053));
NAND2BXL inst_cellmath__24_0_I1835 (.Y(N3346), .AN(N3054), .B(N3055));
NAND2BXL inst_cellmath__24_0_I1838 (.Y(N3349), .AN(N3056), .B(N3057));
NAND2BXL inst_cellmath__24_0_I1841 (.Y(N3352), .AN(N3058), .B(N3059));
NAND2BXL inst_cellmath__24_0_I1844 (.Y(N3355), .AN(N3060), .B(N3061));
NAND2BXL inst_cellmath__24_0_I1847 (.Y(N3358), .AN(N3062), .B(N3063));
NAND2BXL inst_cellmath__24_0_I1850 (.Y(N3361), .AN(N3064), .B(N3065));
NAND2BXL inst_cellmath__24_0_I1853 (.Y(N3364), .AN(N3066), .B(N3067));
NAND2BXL inst_cellmath__24_0_I1856 (.Y(N3367), .AN(N3068), .B(N3069));
NAND2BXL inst_cellmath__24_0_I1859 (.Y(N3370), .AN(N3070), .B(N3071));
NAND2BXL inst_cellmath__24_0_I1862 (.Y(N3373), .AN(N3072), .B(N3073));
NAND2BXL inst_cellmath__24_0_I1865 (.Y(N3376), .AN(N3074), .B(N3075));
NAND2BXL inst_cellmath__24_0_I1868 (.Y(N3379), .AN(N3076), .B(N3077));
NAND2BXL inst_cellmath__24_0_I1871 (.Y(N3382), .AN(N3078), .B(N3079));
NAND2BXL inst_cellmath__24_0_I1874 (.Y(N3385), .AN(N3080), .B(N3081));
NAND2BXL inst_cellmath__24_0_I1877 (.Y(N3388), .AN(N3082), .B(N3083));
NAND2BXL inst_cellmath__24_0_I1880 (.Y(N3391), .AN(N3084), .B(N3085));
NAND2BXL inst_cellmath__24_0_I1883 (.Y(N3394), .AN(N3086), .B(N3087));
NAND2BXL inst_cellmath__24_0_I1886 (.Y(N3397), .AN(N3088), .B(N3089));
NAND2BXL inst_cellmath__24_0_I1889 (.Y(N3400), .AN(N3090), .B(N3091));
NAND2BXL inst_cellmath__24_0_I1892 (.Y(N3403), .AN(N3092), .B(N3093));
NAND2BXL inst_cellmath__24_0_I1895 (.Y(N3406), .AN(N3094), .B(N3095));
NAND2BXL inst_cellmath__24_0_I1898 (.Y(N3409), .AN(N3096), .B(N3097));
NAND2BXL inst_cellmath__24_0_I1901 (.Y(N3412), .AN(N3098), .B(N3099));
NAND2BXL inst_cellmath__24_0_I1904 (.Y(N3415), .AN(N3100), .B(N3101));
NAND2BXL inst_cellmath__24_0_I1907 (.Y(N3418), .AN(N3102), .B(N3103));
NAND2BXL inst_cellmath__24_0_I1910 (.Y(N3421), .AN(N3104), .B(N3105));
NAND2BXL inst_cellmath__24_0_I1913 (.Y(N3424), .AN(N3106), .B(N3107));
NAND2BXL inst_cellmath__24_0_I1916 (.Y(N3427), .AN(N3108), .B(N3109));
XOR2XL inst_cellmath__24_0_I2720 (.Y(inst_cellmath__24_0_out0[15]), .A(N3046), .B(N3337));
XNOR2X1 inst_cellmath__24_0_I1922 (.Y(inst_cellmath__24_0_out0[16]), .A(N4299), .B(N3340));
XNOR2X1 inst_cellmath__24_0_I1923 (.Y(inst_cellmath__24_0_out0[20]), .A(N3246), .B(N3352));
XNOR2X1 inst_cellmath__24_0_I1924 (.Y(inst_cellmath__24_0_out0[22]), .A(N4322), .B(N3358));
XNOR2X1 inst_cellmath__24_0_I1925 (.Y(inst_cellmath__24_0_out0[24]), .A(N4323), .B(N3364));
XNOR2X1 inst_cellmath__24_0_I1926 (.Y(inst_cellmath__24_0_out0[26]), .A(N3284), .B(N3370));
XNOR2X1 inst_cellmath__24_0_I1927 (.Y(inst_cellmath__24_0_out0[28]), .A(N3286), .B(N3376));
XNOR2X1 inst_cellmath__24_0_I1928 (.Y(inst_cellmath__24_0_out0[30]), .A(N3288), .B(N3382));
XNOR2X1 inst_cellmath__24_0_I1929 (.Y(inst_cellmath__24_0_out0[32]), .A(N4325), .B(N3388));
XOR2XL inst_cellmath__24_0_I6148 (.Y(inst_cellmath__24_0_out0[36]), .A(N3326), .B(N3400));
XOR2XL inst_cellmath__24_0_I1931 (.Y(inst_cellmath__24_0_out0[40]), .A(N3328), .B(N3412));
XNOR2X1 inst_cellmath__24_0_I1932 (.Y(inst_cellmath__24_0_out0[44]), .A(N4344), .B(N3424));
XNOR2X1 node_cs_reduced_local_A_I1995 (.Y(N3445), .A(N3343), .B(N3051));
XNOR2X1 node_cs_reduced_local_A_I1996 (.Y(N3446), .A(N3343), .B(N3050));
MXI2XL inst_cellmath__24_0_I1934 (.Y(inst_cellmath__24_0_out0[17]), .A(N3445), .B(N3446), .S0(N4299));
XNOR2X1 node_cs_local_A_I1997 (.Y(N3448), .A(N3346), .B(N4228));
NOR2BX1 node_cs_local_A_I2721 (.Y(N3623), .AN(N3118), .B(N4228));
XOR2XL node_cs_local_A_I1999 (.Y(N3449), .A(N3346), .B(N3623));
MXI2XL inst_cellmath__24_0_I1936 (.Y(inst_cellmath__24_0_out0[18]), .A(N3449), .B(N3448), .S0(N4299));
XNOR2X1 node_cs_local_A_I2000 (.Y(N3451), .A(N3349), .B(N3127));
NOR2XL andori2bb1_A_I2861 (.Y(N4374), .A(N4225), .B(N3118));
NOR2XL andori2bb1_A_I2862 (.Y(N3632), .A(N4374), .B(N3127));
XOR2XL node_cs_local_A_I2002 (.Y(N3452), .A(N3349), .B(N3632));
MXI2XL inst_cellmath__24_0_I1938 (.Y(inst_cellmath__24_0_out0[19]), .A(N3452), .B(N3451), .S0(N4299));
XNOR2X1 node_cs_reduced_local_A_I2003 (.Y(N3454), .A(N3355), .B(N3059));
XNOR2X1 node_cs_reduced_local_A_I2004 (.Y(N3455), .A(N3355), .B(N3058));
MXI2XL inst_cellmath__24_0_I1940 (.Y(inst_cellmath__24_0_out0[21]), .A(N3454), .B(N3455), .S0(N3246));
XNOR2X1 node_cs_reduced_local_A_I2005 (.Y(N3457), .A(N3361), .B(N3063));
XNOR2X1 node_cs_reduced_local_A_I2006 (.Y(N3458), .A(N3361), .B(N3062));
MXI2XL inst_cellmath__24_0_I1942 (.Y(inst_cellmath__24_0_out0[23]), .A(N3457), .B(N3458), .S0(N4322));
XNOR2X1 node_cs_reduced_local_A_I2007 (.Y(N3460), .A(N3367), .B(N3067));
XNOR2X1 node_cs_reduced_local_A_I2722 (.Y(N3461), .A(N3066), .B(N3367));
MXI2XL inst_cellmath__24_0_I1944 (.Y(inst_cellmath__24_0_out0[25]), .A(N3460), .B(N3461), .S0(N4323));
XNOR2X1 node_cs_reduced_local_A_I2009 (.Y(N3463), .A(N3373), .B(N3071));
XNOR2X1 node_cs_reduced_local_A_I2010 (.Y(N3464), .A(N3373), .B(N3070));
MXI2XL inst_cellmath__24_0_I1946 (.Y(inst_cellmath__24_0_out0[27]), .A(N3463), .B(N3464), .S0(N3284));
XNOR2X1 node_cs_reduced_local_A_I2011 (.Y(N3466), .A(N3379), .B(N3075));
XNOR2X1 node_cs_reduced_local_A_I2012 (.Y(N3467), .A(N3379), .B(N3074));
MXI2XL inst_cellmath__24_0_I1948 (.Y(inst_cellmath__24_0_out0[29]), .A(N3466), .B(N3467), .S0(N3286));
XNOR2X1 node_cs_reduced_local_A_I2013 (.Y(N3469), .A(N3385), .B(N3079));
XNOR2X1 node_cs_reduced_local_A_I2014 (.Y(N3470), .A(N3385), .B(N3078));
MXI2XL inst_cellmath__24_0_I1950 (.Y(inst_cellmath__24_0_out0[31]), .A(N3469), .B(N3470), .S0(N3288));
XNOR2X1 node_cs_reduced_local_A_I2015 (.Y(N3472), .A(N3391), .B(N3083));
XNOR2X1 node_cs_reduced_local_A_I2016 (.Y(N3473), .A(N3391), .B(N3082));
MXI2XL inst_cellmath__24_0_I1952 (.Y(inst_cellmath__24_0_out0[33]), .A(N3472), .B(N3473), .S0(N4325));
XNOR2X1 node_cs_local_A_I2017 (.Y(N3475), .A(N3394), .B(N4248));
NOR2BX1 node_cs_local_A_I2723 (.Y(N3690), .AN(N3158), .B(N4248));
XOR2XL node_cs_local_A_I2019 (.Y(N3476), .A(N3394), .B(N3690));
MXI2XL inst_cellmath__24_0_I1954 (.Y(inst_cellmath__24_0_out0[34]), .A(N3476), .B(N3475), .S0(N4325));
XNOR2X1 node_cs_local_A_I2020 (.Y(N3478), .A(N3397), .B(N3167));
NOR2XL andori2bb1_A_I2863 (.Y(N4381), .A(N4245), .B(N3158));
NOR2XL andori2bb1_A_I2864 (.Y(N3699), .A(N4381), .B(N3167));
XOR2XL node_cs_local_A_I2022 (.Y(N3479), .A(N3397), .B(N3699));
MXI2XL inst_cellmath__24_0_I1956 (.Y(inst_cellmath__24_0_out0[35]), .A(N3479), .B(N3478), .S0(N4325));
XNOR2X1 node_cs_reduced_local_A_I2023 (.Y(N3481), .A(N3403), .B(N3091));
XNOR2X1 node_cs_reduced_local_A_I2024 (.Y(N3482), .A(N3403), .B(N3090));
MXI2XL inst_cellmath__24_0_I1958 (.Y(inst_cellmath__24_0_out0[37]), .A(N3482), .B(N3481), .S0(N3326));
XNOR2X1 node_cs_local_A_I2025 (.Y(N3484), .A(N3406), .B(N4256));
NOR2BX1 node_cs_local_A_I2724 (.Y(N3715), .AN(N3174), .B(N4256));
XOR2XL node_cs_local_A_I2027 (.Y(N3485), .A(N3406), .B(N3715));
MXI2XL inst_cellmath__24_0_I1960 (.Y(inst_cellmath__24_0_out0[38]), .A(N3484), .B(N3485), .S0(N3326));
XNOR2X1 node_cs_local_A_I2028 (.Y(N3487), .A(N3409), .B(N3183));
NOR2XL andori2bb1_A_I2865 (.Y(N4388), .A(N4253), .B(N3174));
NOR2XL andori2bb1_A_I2866 (.Y(N3724), .A(N4388), .B(N3183));
XOR2XL node_cs_local_A_I2030 (.Y(N3488), .A(N3409), .B(N3724));
MXI2XL inst_cellmath__24_0_I1962 (.Y(inst_cellmath__24_0_out0[39]), .A(N3487), .B(N3488), .S0(N3326));
XNOR2X1 node_cs_reduced_local_A_I2031 (.Y(N3490), .A(N3415), .B(N3099));
XNOR2X1 node_cs_reduced_local_A_I2032 (.Y(N3491), .A(N3415), .B(N3098));
MXI2XL inst_cellmath__24_0_I1964 (.Y(inst_cellmath__24_0_out0[41]), .A(N3491), .B(N3490), .S0(N3328));
XNOR2X1 node_cs_local_A_I2033 (.Y(N3493), .A(N3418), .B(N4264));
NOR2BX1 node_cs_local_A_I2725 (.Y(N3740), .AN(N3190), .B(N4264));
XOR2XL node_cs_local_A_I2035 (.Y(N3494), .A(N3418), .B(N3740));
MXI2XL inst_cellmath__24_0_I1966 (.Y(inst_cellmath__24_0_out0[42]), .A(N3493), .B(N3494), .S0(N3328));
XNOR2X1 node_cs_local_A_I2036 (.Y(N3496), .A(N3421), .B(N3199));
NOR2XL andori2bb1_A_I2867 (.Y(N4395), .A(N4261), .B(N3190));
NOR2XL andori2bb1_A_I2868 (.Y(N3749), .A(N4395), .B(N3199));
XOR2XL node_cs_local_A_I2038 (.Y(N3497), .A(N3421), .B(N3749));
MXI2XL inst_cellmath__24_0_I1968 (.Y(inst_cellmath__24_0_out0[43]), .A(N3496), .B(N3497), .S0(N3328));
XNOR2X1 node_cs_reduced_local_A_I2039 (.Y(N3499), .A(N3427), .B(N3107));
XNOR2X1 node_cs_reduced_local_A_I2040 (.Y(N3500), .A(N3427), .B(N3106));
MXI2XL inst_cellmath__24_0_I1970 (.Y(inst_cellmath__24_0_out0[45]), .A(N3499), .B(N3500), .S0(N4344));
XNOR2X1 node_cs_local_A_I2041 (.Y(N3502), .A(N3110), .B(N4272));
NOR2BX1 node_cs_local_A_I2726 (.Y(N3765), .AN(N3206), .B(N4272));
XOR2XL node_cs_local_A_I2043 (.Y(N3503), .A(N3110), .B(N3765));
MXI2XL inst_cellmath__24_0_I1972 (.Y(inst_cellmath__24_0_out0[46]), .A(N3503), .B(N3502), .S0(N4344));
AOI21X4 inst_cellmath__24_0_I1992 (.Y(inst_cellmath__24_0_out0[47]), .A0(N3215), .A1(N3330), .B0(N3505));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw3815070899_bdw (
	inst_cellmath__25_0_out0,
	inst_cellmath__25_0_in0
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__25_0_out0;
input [47:0] inst_cellmath__25_0_in0;
wire N146,N147,N148,N149,N150,N151,N152 
	,N153,N154,N155,N156,N157,N158,N159,N160 
	,N161,N162,N163,N164,N165,N166,N167,N168 
	,N169,N170,N171,N172,N173,N174,N175,N176 
	,N177,N178,N179,N180,N181,N182,N183,N184 
	,N185,N186,N187,N188,N189,N190,N191,N192 
	,N294,N297,N298,N299,N300,N301,N302;
INVXL inst_cellmath__25_0_I0 (.Y(N146), .A(inst_cellmath__25_0_in0[0]));
INVXL inst_cellmath__25_0_I1 (.Y(N147), .A(inst_cellmath__25_0_in0[1]));
INVXL inst_cellmath__25_0_I2 (.Y(N148), .A(inst_cellmath__25_0_in0[2]));
INVXL inst_cellmath__25_0_I3 (.Y(N149), .A(inst_cellmath__25_0_in0[3]));
INVXL inst_cellmath__25_0_I4 (.Y(N150), .A(inst_cellmath__25_0_in0[4]));
INVXL inst_cellmath__25_0_I5 (.Y(N151), .A(inst_cellmath__25_0_in0[5]));
INVXL inst_cellmath__25_0_I6 (.Y(N152), .A(inst_cellmath__25_0_in0[6]));
INVXL inst_cellmath__25_0_I7 (.Y(N153), .A(inst_cellmath__25_0_in0[7]));
INVXL inst_cellmath__25_0_I8 (.Y(N154), .A(inst_cellmath__25_0_in0[8]));
INVXL inst_cellmath__25_0_I9 (.Y(N155), .A(inst_cellmath__25_0_in0[9]));
INVXL inst_cellmath__25_0_I10 (.Y(N156), .A(inst_cellmath__25_0_in0[10]));
INVXL inst_cellmath__25_0_I11 (.Y(N157), .A(inst_cellmath__25_0_in0[11]));
INVXL inst_cellmath__25_0_I12 (.Y(N158), .A(inst_cellmath__25_0_in0[12]));
INVXL inst_cellmath__25_0_I13 (.Y(N159), .A(inst_cellmath__25_0_in0[13]));
INVXL inst_cellmath__25_0_I14 (.Y(N160), .A(inst_cellmath__25_0_in0[14]));
INVXL inst_cellmath__25_0_I15 (.Y(N161), .A(inst_cellmath__25_0_in0[15]));
INVXL inst_cellmath__25_0_I16 (.Y(N162), .A(inst_cellmath__25_0_in0[16]));
INVXL inst_cellmath__25_0_I17 (.Y(N163), .A(inst_cellmath__25_0_in0[17]));
INVXL inst_cellmath__25_0_I18 (.Y(N164), .A(inst_cellmath__25_0_in0[18]));
INVXL inst_cellmath__25_0_I19 (.Y(N165), .A(inst_cellmath__25_0_in0[19]));
INVXL inst_cellmath__25_0_I20 (.Y(N166), .A(inst_cellmath__25_0_in0[20]));
INVXL inst_cellmath__25_0_I21 (.Y(N167), .A(inst_cellmath__25_0_in0[21]));
INVXL inst_cellmath__25_0_I22 (.Y(N168), .A(inst_cellmath__25_0_in0[22]));
INVXL inst_cellmath__25_0_I23 (.Y(N169), .A(inst_cellmath__25_0_in0[23]));
INVXL inst_cellmath__25_0_I24 (.Y(N170), .A(inst_cellmath__25_0_in0[24]));
INVXL inst_cellmath__25_0_I25 (.Y(N171), .A(inst_cellmath__25_0_in0[25]));
INVXL inst_cellmath__25_0_I26 (.Y(N172), .A(inst_cellmath__25_0_in0[26]));
INVXL inst_cellmath__25_0_I27 (.Y(N173), .A(inst_cellmath__25_0_in0[27]));
INVXL inst_cellmath__25_0_I28 (.Y(N174), .A(inst_cellmath__25_0_in0[28]));
INVXL inst_cellmath__25_0_I29 (.Y(N175), .A(inst_cellmath__25_0_in0[29]));
INVXL inst_cellmath__25_0_I30 (.Y(N176), .A(inst_cellmath__25_0_in0[30]));
INVXL inst_cellmath__25_0_I31 (.Y(N177), .A(inst_cellmath__25_0_in0[31]));
INVXL inst_cellmath__25_0_I32 (.Y(N178), .A(inst_cellmath__25_0_in0[32]));
INVXL inst_cellmath__25_0_I33 (.Y(N179), .A(inst_cellmath__25_0_in0[33]));
INVXL inst_cellmath__25_0_I34 (.Y(N180), .A(inst_cellmath__25_0_in0[34]));
INVXL inst_cellmath__25_0_I35 (.Y(N181), .A(inst_cellmath__25_0_in0[35]));
INVXL inst_cellmath__25_0_I36 (.Y(N182), .A(inst_cellmath__25_0_in0[36]));
INVXL inst_cellmath__25_0_I37 (.Y(N183), .A(inst_cellmath__25_0_in0[37]));
INVXL inst_cellmath__25_0_I38 (.Y(N184), .A(inst_cellmath__25_0_in0[38]));
INVXL inst_cellmath__25_0_I39 (.Y(N185), .A(inst_cellmath__25_0_in0[39]));
INVXL inst_cellmath__25_0_I40 (.Y(N186), .A(inst_cellmath__25_0_in0[40]));
INVXL inst_cellmath__25_0_I41 (.Y(N187), .A(inst_cellmath__25_0_in0[41]));
INVXL inst_cellmath__25_0_I42 (.Y(N188), .A(inst_cellmath__25_0_in0[42]));
INVXL inst_cellmath__25_0_I43 (.Y(N189), .A(inst_cellmath__25_0_in0[43]));
INVXL inst_cellmath__25_0_I44 (.Y(N190), .A(inst_cellmath__25_0_in0[44]));
INVXL inst_cellmath__25_0_I45 (.Y(N191), .A(inst_cellmath__25_0_in0[45]));
INVXL inst_cellmath__25_0_I46 (.Y(N192), .A(inst_cellmath__25_0_in0[46]));
CLKINVX6 inst_cellmath__25_0_I145 (.Y(N294), .A(inst_cellmath__25_0_in0[47]));
INVX2 inst_cellmath__25_0_I153 (.Y(N302), .A(N294));
NOR2BX1 inst_cellmath__25_0_I96 (.Y(inst_cellmath__25_0_out0[0]), .AN(N302), .B(N146));
MXI2XL inst_cellmath__25_0_I97 (.Y(inst_cellmath__25_0_out0[1]), .A(N146), .B(N147), .S0(N302));
MXI2XL inst_cellmath__25_0_I98 (.Y(inst_cellmath__25_0_out0[2]), .A(N147), .B(N148), .S0(N302));
MXI2XL inst_cellmath__25_0_I99 (.Y(inst_cellmath__25_0_out0[3]), .A(N148), .B(N149), .S0(N302));
MXI2XL inst_cellmath__25_0_I100 (.Y(inst_cellmath__25_0_out0[4]), .A(N149), .B(N150), .S0(N302));
INVX2 inst_cellmath__25_0_I152 (.Y(N301), .A(N294));
MXI2XL inst_cellmath__25_0_I101 (.Y(inst_cellmath__25_0_out0[5]), .A(N150), .B(N151), .S0(N301));
MXI2XL inst_cellmath__25_0_I102 (.Y(inst_cellmath__25_0_out0[6]), .A(N151), .B(N152), .S0(N301));
MXI2XL inst_cellmath__25_0_I103 (.Y(inst_cellmath__25_0_out0[7]), .A(N152), .B(N153), .S0(N301));
MXI2XL inst_cellmath__25_0_I104 (.Y(inst_cellmath__25_0_out0[8]), .A(N153), .B(N154), .S0(N301));
MXI2XL inst_cellmath__25_0_I105 (.Y(inst_cellmath__25_0_out0[9]), .A(N154), .B(N155), .S0(N301));
MXI2XL inst_cellmath__25_0_I106 (.Y(inst_cellmath__25_0_out0[10]), .A(N155), .B(N156), .S0(N301));
INVX3 inst_cellmath__25_0_I151 (.Y(N300), .A(N294));
MXI2XL inst_cellmath__25_0_I107 (.Y(inst_cellmath__25_0_out0[11]), .A(N156), .B(N157), .S0(N300));
MXI2XL inst_cellmath__25_0_I108 (.Y(inst_cellmath__25_0_out0[12]), .A(N157), .B(N158), .S0(N300));
MXI2XL inst_cellmath__25_0_I109 (.Y(inst_cellmath__25_0_out0[13]), .A(N158), .B(N159), .S0(N300));
MXI2XL inst_cellmath__25_0_I110 (.Y(inst_cellmath__25_0_out0[14]), .A(N159), .B(N160), .S0(N300));
MXI2XL inst_cellmath__25_0_I111 (.Y(inst_cellmath__25_0_out0[15]), .A(N160), .B(N161), .S0(N300));
MXI2X1 inst_cellmath__25_0_I112 (.Y(inst_cellmath__25_0_out0[16]), .A(N161), .B(N162), .S0(N300));
CLKINVX4 inst_cellmath__25_0_I150 (.Y(N299), .A(N294));
MXI2XL inst_cellmath__25_0_I113 (.Y(inst_cellmath__25_0_out0[17]), .A(N162), .B(N163), .S0(N299));
MXI2X1 inst_cellmath__25_0_I114 (.Y(inst_cellmath__25_0_out0[18]), .A(N163), .B(N164), .S0(N299));
MXI2XL inst_cellmath__25_0_I115 (.Y(inst_cellmath__25_0_out0[19]), .A(N164), .B(N165), .S0(N299));
MXI2XL inst_cellmath__25_0_I116 (.Y(inst_cellmath__25_0_out0[20]), .A(N165), .B(N166), .S0(N299));
MXI2XL inst_cellmath__25_0_I117 (.Y(inst_cellmath__25_0_out0[21]), .A(N166), .B(N167), .S0(N299));
MXI2X1 inst_cellmath__25_0_I118 (.Y(inst_cellmath__25_0_out0[22]), .A(N167), .B(N168), .S0(N299));
INVXL inst_cellmath__25_0_I149 (.Y(N298), .A(N294));
MXI2XL inst_cellmath__25_0_I119 (.Y(inst_cellmath__25_0_out0[23]), .A(N168), .B(N169), .S0(N298));
MXI2X1 inst_cellmath__25_0_I120 (.Y(inst_cellmath__25_0_out0[24]), .A(N169), .B(N170), .S0(N298));
MXI2XL inst_cellmath__25_0_I121 (.Y(inst_cellmath__25_0_out0[25]), .A(N170), .B(N171), .S0(N298));
MXI2XL inst_cellmath__25_0_I122 (.Y(inst_cellmath__25_0_out0[26]), .A(N171), .B(N172), .S0(N298));
MXI2XL inst_cellmath__25_0_I123 (.Y(inst_cellmath__25_0_out0[27]), .A(N172), .B(N173), .S0(N298));
MXI2XL inst_cellmath__25_0_I124 (.Y(inst_cellmath__25_0_out0[28]), .A(N173), .B(N174), .S0(N298));
INVXL inst_cellmath__25_0_I148 (.Y(N297), .A(N294));
MXI2XL inst_cellmath__25_0_I125 (.Y(inst_cellmath__25_0_out0[29]), .A(N174), .B(N175), .S0(N297));
MXI2XL inst_cellmath__25_0_I126 (.Y(inst_cellmath__25_0_out0[30]), .A(N175), .B(N176), .S0(N297));
MXI2XL inst_cellmath__25_0_I127 (.Y(inst_cellmath__25_0_out0[31]), .A(N176), .B(N177), .S0(N297));
MXI2XL inst_cellmath__25_0_I128 (.Y(inst_cellmath__25_0_out0[32]), .A(N177), .B(N178), .S0(N297));
MXI2XL inst_cellmath__25_0_I129 (.Y(inst_cellmath__25_0_out0[33]), .A(N178), .B(N179), .S0(N297));
MXI2XL inst_cellmath__25_0_I130 (.Y(inst_cellmath__25_0_out0[34]), .A(N179), .B(N180), .S0(N297));
MXI2XL inst_cellmath__25_0_I131 (.Y(inst_cellmath__25_0_out0[35]), .A(N180), .B(N181), .S0(N297));
MXI2XL inst_cellmath__25_0_I132 (.Y(inst_cellmath__25_0_out0[36]), .A(N181), .B(N182), .S0(N297));
MXI2XL inst_cellmath__25_0_I133 (.Y(inst_cellmath__25_0_out0[37]), .A(N182), .B(N183), .S0(N297));
MXI2XL inst_cellmath__25_0_I134 (.Y(inst_cellmath__25_0_out0[38]), .A(N183), .B(N184), .S0(N297));
MXI2XL inst_cellmath__25_0_I135 (.Y(inst_cellmath__25_0_out0[39]), .A(N184), .B(N185), .S0(N297));
MXI2XL inst_cellmath__25_0_I136 (.Y(inst_cellmath__25_0_out0[40]), .A(N185), .B(N186), .S0(N297));
MXI2XL inst_cellmath__25_0_I137 (.Y(inst_cellmath__25_0_out0[41]), .A(N186), .B(N187), .S0(N298));
MXI2XL inst_cellmath__25_0_I138 (.Y(inst_cellmath__25_0_out0[42]), .A(N187), .B(N188), .S0(N298));
MXI2XL inst_cellmath__25_0_I139 (.Y(inst_cellmath__25_0_out0[43]), .A(N188), .B(N189), .S0(N298));
MXI2XL inst_cellmath__25_0_I140 (.Y(inst_cellmath__25_0_out0[44]), .A(N189), .B(N190), .S0(N298));
MXI2XL inst_cellmath__25_0_I141 (.Y(inst_cellmath__25_0_out0[45]), .A(N190), .B(N191), .S0(N298));
MXI2XL inst_cellmath__25_0_I142 (.Y(inst_cellmath__25_0_out0[46]), .A(N191), .B(N192), .S0(N298));
NAND2BXL inst_cellmath__25_0_I154 (.Y(inst_cellmath__25_0_out0[47]), .AN(N302), .B(N192));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw3815070899_bdw (
	inst_cellmath__45_0_out0,
	inst_cellmath__45_0_in0
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__45_0_out0;
input [47:24] inst_cellmath__45_0_in0;
wire N150,N152,N154,N156,N158,N160,N162 
	,N164,N166,N168,N170,N172,N174,N176,N178 
	,N180,N182,N184,N186,N188,N192,N197,N201 
	,N208,N210,N212,N214,N216,N218,N220,N222 
	,N224,N226,N228,N230,N232,N234,N236,N238 
	,N242,N246,N255,N259,N262,N265,N272,N274 
	,N276,N278,N280,N282,N284,N286,N294,N300 
	,N302,N319,N323,N356,N395,N399,N402,N405 
	,N408,N414,N417,N738,N739,N740,N745,N748 
	,N749,N750,N751,N754,N755,N756,N757,N758 
	,N817,N823,N830,N837,N844;
AND2XL inst_cellmath__45_0_I39 (.Y(N197), .A(inst_cellmath__45_0_in0[25]), .B(inst_cellmath__45_0_in0[24]));
AND2XL inst_cellmath__45_0_I42 (.Y(N150), .A(inst_cellmath__45_0_in0[26]), .B(inst_cellmath__45_0_in0[25]));
AND2XL inst_cellmath__45_0_I44 (.Y(N152), .A(inst_cellmath__45_0_in0[27]), .B(inst_cellmath__45_0_in0[26]));
AND2XL inst_cellmath__45_0_I46 (.Y(N154), .A(inst_cellmath__45_0_in0[28]), .B(inst_cellmath__45_0_in0[27]));
AND2XL inst_cellmath__45_0_I48 (.Y(N156), .A(inst_cellmath__45_0_in0[29]), .B(inst_cellmath__45_0_in0[28]));
AND2XL inst_cellmath__45_0_I50 (.Y(N158), .A(inst_cellmath__45_0_in0[30]), .B(inst_cellmath__45_0_in0[29]));
AND2XL inst_cellmath__45_0_I52 (.Y(N160), .A(inst_cellmath__45_0_in0[31]), .B(inst_cellmath__45_0_in0[30]));
AND2XL inst_cellmath__45_0_I54 (.Y(N162), .A(inst_cellmath__45_0_in0[32]), .B(inst_cellmath__45_0_in0[31]));
AND2XL inst_cellmath__45_0_I56 (.Y(N164), .A(inst_cellmath__45_0_in0[33]), .B(inst_cellmath__45_0_in0[32]));
AND2XL inst_cellmath__45_0_I58 (.Y(N166), .A(inst_cellmath__45_0_in0[34]), .B(inst_cellmath__45_0_in0[33]));
AND2XL inst_cellmath__45_0_I60 (.Y(N168), .A(inst_cellmath__45_0_in0[35]), .B(inst_cellmath__45_0_in0[34]));
AND2XL inst_cellmath__45_0_I62 (.Y(N170), .A(inst_cellmath__45_0_in0[36]), .B(inst_cellmath__45_0_in0[35]));
CLKAND2X2 inst_cellmath__45_0_I64 (.Y(N172), .A(inst_cellmath__45_0_in0[37]), .B(inst_cellmath__45_0_in0[36]));
AND2XL inst_cellmath__45_0_I66 (.Y(N174), .A(inst_cellmath__45_0_in0[38]), .B(inst_cellmath__45_0_in0[37]));
AND2XL inst_cellmath__45_0_I68 (.Y(N176), .A(inst_cellmath__45_0_in0[39]), .B(inst_cellmath__45_0_in0[38]));
AND2XL inst_cellmath__45_0_I70 (.Y(N178), .A(inst_cellmath__45_0_in0[40]), .B(inst_cellmath__45_0_in0[39]));
CLKAND2X2 inst_cellmath__45_0_I72 (.Y(N180), .A(inst_cellmath__45_0_in0[41]), .B(inst_cellmath__45_0_in0[40]));
AND2XL inst_cellmath__45_0_I74 (.Y(N182), .A(inst_cellmath__45_0_in0[42]), .B(inst_cellmath__45_0_in0[41]));
AND2X1 inst_cellmath__45_0_I76 (.Y(N184), .A(inst_cellmath__45_0_in0[42]), .B(inst_cellmath__45_0_in0[43]));
AND2XL inst_cellmath__45_0_I78 (.Y(N186), .A(inst_cellmath__45_0_in0[44]), .B(inst_cellmath__45_0_in0[43]));
AND2XL inst_cellmath__45_0_I80 (.Y(N188), .A(inst_cellmath__45_0_in0[45]), .B(inst_cellmath__45_0_in0[44]));
AND2XL inst_cellmath__45_0_I84 (.Y(N192), .A(inst_cellmath__45_0_in0[47]), .B(inst_cellmath__45_0_in0[46]));
INVXL inst_cellmath__45_0_I412 (.Y(inst_cellmath__45_0_out0[0]), .A(inst_cellmath__45_0_in0[24]));
NAND2XL inst_cellmath__45_0_I91 (.Y(N201), .A(N150), .B(inst_cellmath__45_0_in0[24]));
AND2XL inst_cellmath__45_0_I93 (.Y(N255), .A(N152), .B(N197));
NAND2XL inst_cellmath__45_0_I96 (.Y(N208), .A(N154), .B(N150));
AND2XL inst_cellmath__45_0_I98 (.Y(N210), .A(N156), .B(N152));
NAND2XL inst_cellmath__45_0_I100 (.Y(N212), .A(N158), .B(N154));
AND2XL inst_cellmath__45_0_I102 (.Y(N214), .A(N160), .B(N156));
NAND2XL inst_cellmath__45_0_I104 (.Y(N216), .A(N162), .B(N158));
AND2XL inst_cellmath__45_0_I106 (.Y(N218), .A(N164), .B(N160));
NAND2XL inst_cellmath__45_0_I108 (.Y(N220), .A(N166), .B(N162));
AND2XL inst_cellmath__45_0_I110 (.Y(N222), .A(N168), .B(N164));
NAND2XL inst_cellmath__45_0_I112 (.Y(N224), .A(N170), .B(N166));
AND2XL inst_cellmath__45_0_I114 (.Y(N226), .A(N172), .B(N168));
NAND2XL inst_cellmath__45_0_I116 (.Y(N228), .A(N174), .B(N170));
CLKAND2X6 inst_cellmath__45_0_I118 (.Y(N230), .A(N176), .B(N172));
NAND2XL inst_cellmath__45_0_I120 (.Y(N232), .A(N178), .B(N174));
AND2XL inst_cellmath__45_0_I122 (.Y(N234), .A(N180), .B(N176));
NAND2XL inst_cellmath__45_0_I124 (.Y(N236), .A(N182), .B(N178));
CLKAND2X6 inst_cellmath__45_0_I126 (.Y(N238), .A(N184), .B(N180));
AND2XL inst_cellmath__45_0_I130 (.Y(N242), .A(N188), .B(N184));
CLKAND2X2 inst_cellmath__45_0_I134 (.Y(N246), .A(N192), .B(N188));
INVXL inst_cellmath__45_0_I415 (.Y(N738), .A(inst_cellmath__45_0_out0[0]));
INVXL inst_cellmath__45_0_I416 (.Y(N739), .A(N197));
INVXL inst_cellmath__45_0_I417 (.Y(N740), .A(N201));
NOR2XL inst_cellmath__45_0_I145 (.Y(N259), .A(N208), .B(inst_cellmath__45_0_out0[0]));
NAND2XL inst_cellmath__45_0_I147 (.Y(N262), .A(N210), .B(N197));
NOR2XL inst_cellmath__45_0_I149 (.Y(N265), .A(N212), .B(N201));
NAND2X1 inst_cellmath__45_0_I151 (.Y(N319), .A(N214), .B(N255));
NOR2XL inst_cellmath__45_0_I154 (.Y(N272), .A(N216), .B(N208));
NAND2XL inst_cellmath__45_0_I156 (.Y(N274), .A(N218), .B(N210));
NOR2XL inst_cellmath__45_0_I158 (.Y(N276), .A(N220), .B(N212));
AND2XL inst_cellmath__45_0_I160 (.Y(N278), .A(N222), .B(N214));
NOR2XL inst_cellmath__45_0_I162 (.Y(N280), .A(N224), .B(N216));
NAND2XL inst_cellmath__45_0_I164 (.Y(N282), .A(N226), .B(N218));
NOR2XL inst_cellmath__45_0_I166 (.Y(N284), .A(N228), .B(N220));
NAND2X8 inst_cellmath__45_0_I168 (.Y(N286), .A(N230), .B(N222));
AND2XL inst_cellmath__45_0_I176 (.Y(N294), .A(N238), .B(N230));
NAND3XL hyperpropagate_4_1_A_I570 (.Y(N817), .A(inst_cellmath__45_0_in0[46]), .B(inst_cellmath__45_0_in0[45]), .C(N186));
NOR2XL hyperpropagate_4_1_A_I571 (.Y(N300), .A(N236), .B(N817));
NAND2X6 inst_cellmath__45_0_I184 (.Y(N302), .A(N246), .B(N238));
INVXL inst_cellmath__45_0_I422 (.Y(N745), .A(N739));
INVXL inst_cellmath__45_0_I425 (.Y(N748), .A(N255));
INVXL inst_cellmath__45_0_I426 (.Y(N749), .A(N259));
INVXL inst_cellmath__45_0_I427 (.Y(N750), .A(N262));
INVXL inst_cellmath__45_0_I428 (.Y(N751), .A(N265));
NAND2XL inst_cellmath__45_0_I203 (.Y(N323), .A(N272), .B(N738));
NOR2XL inst_cellmath__45_0_I501 (.Y(N395), .A(N286), .B(N319));
NAND4BXL inst_cellmath__45_0_I506 (.Y(N356), .AN(N232), .B(N186), .C(N280), .D(N182));
AND2XL inst_cellmath__45_0_I509 (.Y(N754), .A(N276), .B(N740));
AND2XL inst_cellmath__45_0_I510 (.Y(N755), .A(N278), .B(N255));
AND2XL inst_cellmath__45_0_I511 (.Y(N756), .A(N280), .B(N259));
OR2XL inst_cellmath__45_0_I512 (.Y(N757), .A(N282), .B(N262));
AND2XL inst_cellmath__45_0_I513 (.Y(N758), .A(N284), .B(N265));
NAND4BBXL inst_cellmath__45_0_I514 (.Y(N399), .AN(N232), .BN(N224), .C(N738), .D(N272));
NAND4BXL inst_cellmath__45_0_I515 (.Y(N402), .AN(N274), .B(N234), .C(N745), .D(N226));
NAND4BBXL inst_cellmath__45_0_I516 (.Y(N405), .AN(N236), .BN(N228), .C(N740), .D(N276));
NAND2XL hyperpropagate_3_1_A_I572 (.Y(N823), .A(N294), .B(N278));
NOR2XL hyperpropagate_3_1_A_I573 (.Y(N408), .A(N748), .B(N823));
NAND4BXL inst_cellmath__45_0_I518 (.Y(N414), .AN(N282), .B(N242), .C(N750), .D(N234));
NAND2XL hyperpropagate_3_1_A_I574 (.Y(N830), .A(N300), .B(N284));
NOR2XL hyperpropagate_3_1_A_I575 (.Y(N417), .A(N751), .B(N830));
NOR3X4 inst_cellmath__45_0_I586 (.Y(inst_cellmath__45_0_out0[24]), .A(N302), .B(N286), .C(N319));
XOR2XL inst_cellmath__45_0_I521 (.Y(inst_cellmath__45_0_out0[1]), .A(N738), .B(inst_cellmath__45_0_in0[25]));
XOR2XL inst_cellmath__45_0_I522 (.Y(inst_cellmath__45_0_out0[2]), .A(N745), .B(inst_cellmath__45_0_in0[26]));
XOR2XL inst_cellmath__45_0_I523 (.Y(inst_cellmath__45_0_out0[3]), .A(N740), .B(inst_cellmath__45_0_in0[27]));
XNOR2X1 inst_cellmath__45_0_I546 (.Y(inst_cellmath__45_0_out0[4]), .A(N748), .B(inst_cellmath__45_0_in0[28]));
XNOR2X1 inst_cellmath__45_0_I364 (.Y(inst_cellmath__45_0_out0[5]), .A(N749), .B(inst_cellmath__45_0_in0[29]));
XOR2XL inst_cellmath__45_0_I525 (.Y(inst_cellmath__45_0_out0[6]), .A(N750), .B(inst_cellmath__45_0_in0[30]));
XNOR2X1 inst_cellmath__45_0_I366 (.Y(inst_cellmath__45_0_out0[7]), .A(N751), .B(inst_cellmath__45_0_in0[31]));
XNOR2X1 inst_cellmath__45_0_I367 (.Y(inst_cellmath__45_0_out0[8]), .A(N319), .B(inst_cellmath__45_0_in0[32]));
XNOR2X1 inst_cellmath__45_0_I368 (.Y(inst_cellmath__45_0_out0[9]), .A(N323), .B(inst_cellmath__45_0_in0[33]));
NOR2XL node_cs_const1_cs_A_I576 (.Y(N837), .A(N274), .B(N739));
XOR2XL node_cs_const1_cs_A_I822 (.Y(inst_cellmath__45_0_out0[10]), .A(inst_cellmath__45_0_in0[34]), .B(N837));
XOR2XL inst_cellmath__45_0_I562 (.Y(inst_cellmath__45_0_out0[11]), .A(N754), .B(inst_cellmath__45_0_in0[35]));
XOR2XL inst_cellmath__45_0_I528 (.Y(inst_cellmath__45_0_out0[12]), .A(N755), .B(inst_cellmath__45_0_in0[36]));
XOR2XL inst_cellmath__45_0_I529 (.Y(inst_cellmath__45_0_out0[13]), .A(N756), .B(inst_cellmath__45_0_in0[37]));
XNOR2X1 inst_cellmath__45_0_I373 (.Y(inst_cellmath__45_0_out0[14]), .A(N757), .B(inst_cellmath__45_0_in0[38]));
XOR2XL inst_cellmath__45_0_I823 (.Y(inst_cellmath__45_0_out0[15]), .A(N758), .B(inst_cellmath__45_0_in0[39]));
XOR2XL inst_cellmath__45_0_I531 (.Y(inst_cellmath__45_0_out0[16]), .A(N395), .B(inst_cellmath__45_0_in0[40]));
XNOR2X1 inst_cellmath__45_0_I376 (.Y(inst_cellmath__45_0_out0[17]), .A(N399), .B(inst_cellmath__45_0_in0[41]));
XNOR2X1 inst_cellmath__45_0_I377 (.Y(inst_cellmath__45_0_out0[18]), .A(N402), .B(inst_cellmath__45_0_in0[42]));
XNOR2X1 inst_cellmath__45_0_I378 (.Y(inst_cellmath__45_0_out0[19]), .A(N405), .B(inst_cellmath__45_0_in0[43]));
XOR2XL inst_cellmath__45_0_I532 (.Y(inst_cellmath__45_0_out0[20]), .A(N408), .B(inst_cellmath__45_0_in0[44]));
NOR2XL node_cs_const1_cs_A_I578 (.Y(N844), .A(N356), .B(N749));
XOR2XL node_cs_const1_cs_A_I824 (.Y(inst_cellmath__45_0_out0[21]), .A(inst_cellmath__45_0_in0[45]), .B(N844));
XNOR2X1 inst_cellmath__45_0_I381 (.Y(inst_cellmath__45_0_out0[22]), .A(N414), .B(inst_cellmath__45_0_in0[46]));
XOR2XL inst_cellmath__45_0_I534 (.Y(inst_cellmath__45_0_out0[23]), .A(N417), .B(inst_cellmath__45_0_in0[47]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw3815070899_bdw (
	inst_cellmath__5_1_out0,
	inst_cellmath__5_1_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__5_1_out0;
input [2:0] inst_cellmath__5_1_in0;
wire N24,N26,N28;
INVXL inst_cellmath__5_1_I11 (.Y(N24), .A(inst_cellmath__5_1_in0[1]));
INVX1 inst_cellmath__5_1_I12 (.Y(N26), .A(inst_cellmath__5_1_in0[2]));
NAND3X1 inst_cellmath__5_1_I13 (.Y(N28), .A(inst_cellmath__5_1_in0[0]), .B(N26), .C(N24));
INVXL inst_cellmath__5_1_I14 (.Y(inst_cellmath__5_1_out0), .A(N28));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw3815070899_bdw (
	inst_cellmath__44__31__out0,
	inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__31__out0;
input  inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1;
wire N13;
INVXL inst_cellmath__44__31__I3 (.Y(N13), .A(inst_cellmath__44__31__in1));
CLKAND2X3 inst_cellmath__44__31__I1 (.Y(inst_cellmath__44__31__out0[0]), .A(inst_cellmath__44__31__in0), .B(N13));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw3815070899_bdw (
	inst_cellmath__6_0_out0,
	inst_cellmath__6_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__6_0_out0;
input [2:0] inst_cellmath__6_0_in0;
wire N29,N34,N36;
INVXL inst_cellmath__6_0_I16 (.Y(N29), .A(inst_cellmath__6_0_in0[0]));
INVX1 inst_cellmath__6_0_I18 (.Y(N34), .A(inst_cellmath__6_0_in0[2]));
NAND3X1 inst_cellmath__6_0_I19 (.Y(N36), .A(inst_cellmath__6_0_in0[1]), .B(N34), .C(N29));
INVXL inst_cellmath__6_0_I20 (.Y(inst_cellmath__6_0_out0), .A(N36));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw3815070899_bdw (
	inst_cellmath__44__30__out0,
	inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__30__out0;
input  inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1;
AND2XL inst_cellmath__44__30__I0 (.Y(inst_cellmath__44__30__out0[0]), .A(inst_cellmath__44__30__in0), .B(inst_cellmath__44__30__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw3815070899_bdw (
	inst_cellmath__8_0_out0,
	inst_cellmath__8_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__8_0_out0;
input [2:0] inst_cellmath__8_0_in0;
wire N30,N32,N37;
INVXL inst_cellmath__8_0_I17 (.Y(N30), .A(inst_cellmath__8_0_in0[0]));
INVX1 inst_cellmath__8_0_I18 (.Y(N32), .A(inst_cellmath__8_0_in0[1]));
NAND3X1 inst_cellmath__8_0_I20 (.Y(N37), .A(inst_cellmath__8_0_in0[2]), .B(N32), .C(N30));
INVXL inst_cellmath__8_0_I21 (.Y(inst_cellmath__8_0_out0), .A(N37));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw3815070899_bdw (
	inst_cellmath__4_0_out0,
	inst_cellmath__4_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__4_0_out0;
input [2:0] inst_cellmath__4_0_in0;
wire N31,N33,N35,N37;
INVX1 inst_cellmath__4_0_I18 (.Y(N31), .A(inst_cellmath__4_0_in0[0]));
CLKINVX1 inst_cellmath__4_0_I19 (.Y(N33), .A(inst_cellmath__4_0_in0[1]));
INVXL inst_cellmath__4_0_I20 (.Y(N35), .A(inst_cellmath__4_0_in0[2]));
NAND3X2 inst_cellmath__4_0_I21 (.Y(N37), .A(N31), .B(N33), .C(N35));
INVX1 inst_cellmath__4_0_I22 (.Y(inst_cellmath__4_0_out0), .A(N37));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw3815070899_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__34_0_out0;
input [22:0] inst_cellmath__34_0_in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48,N49 
	;
NOR2X1 inst_cellmath__34_0_I0 (.Y(N26), .A(inst_cellmath__34_0_in0[0]), .B(inst_cellmath__34_0_in0[1]));
NOR2X1 inst_cellmath__34_0_I1 (.Y(N27), .A(inst_cellmath__34_0_in0[22]), .B(inst_cellmath__34_0_in0[21]));
NOR2X1 inst_cellmath__34_0_I2 (.Y(N28), .A(inst_cellmath__34_0_in0[20]), .B(inst_cellmath__34_0_in0[19]));
NOR2X2 inst_cellmath__34_0_I3 (.Y(N29), .A(inst_cellmath__34_0_in0[18]), .B(inst_cellmath__34_0_in0[17]));
NOR2X2 inst_cellmath__34_0_I4 (.Y(N30), .A(inst_cellmath__34_0_in0[16]), .B(inst_cellmath__34_0_in0[15]));
NOR2X1 inst_cellmath__34_0_I5 (.Y(N31), .A(inst_cellmath__34_0_in0[14]), .B(inst_cellmath__34_0_in0[13]));
NOR2X1 inst_cellmath__34_0_I6 (.Y(N32), .A(inst_cellmath__34_0_in0[12]), .B(inst_cellmath__34_0_in0[11]));
NOR2XL inst_cellmath__34_0_I7 (.Y(N33), .A(inst_cellmath__34_0_in0[10]), .B(inst_cellmath__34_0_in0[9]));
NOR2XL inst_cellmath__34_0_I8 (.Y(N34), .A(inst_cellmath__34_0_in0[8]), .B(inst_cellmath__34_0_in0[7]));
NOR2XL inst_cellmath__34_0_I9 (.Y(N35), .A(inst_cellmath__34_0_in0[6]), .B(inst_cellmath__34_0_in0[5]));
NOR2XL inst_cellmath__34_0_I10 (.Y(N36), .A(inst_cellmath__34_0_in0[4]), .B(inst_cellmath__34_0_in0[3]));
INVXL inst_cellmath__34_0_I11 (.Y(N37), .A(inst_cellmath__34_0_in0[2]));
NAND2X2 inst_cellmath__34_0_I12 (.Y(N38), .A(N37), .B(N26));
NAND2X2 inst_cellmath__34_0_I13 (.Y(N39), .A(N27), .B(N28));
NAND2X4 inst_cellmath__34_0_I14 (.Y(N40), .A(N29), .B(N30));
NAND2X2 inst_cellmath__34_0_I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__34_0_I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__34_0_I17 (.Y(N43), .A(N35), .B(N36));
NOR2X2 inst_cellmath__34_0_I18 (.Y(N44), .A(N38), .B(N39));
NOR2X4 inst_cellmath__34_0_I19 (.Y(N45), .A(N40), .B(N41));
NAND2X2 inst_cellmath__34_0_I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__34_0_I180 (.Y(N48), .A(N42), .B(N43));
NOR2X2 inst_cellmath__34_0_I23 (.Y(N49), .A(N48), .B(N47));
INVX2 inst_cellmath__34_0_I24 (.Y(inst_cellmath__34_0_out0), .A(N49));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw3815070899_bdw (
	inst_cellmath__44__29__out0,
	inst_cellmath__44__29__in0,
	inst_cellmath__44__29__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__29__out0;
input  inst_cellmath__44__29__in0;
input [24:24] inst_cellmath__44__29__in1;
wire N5;
NOR2X2 inst_cellmath__44__29__I0 (.Y(N5), .A(inst_cellmath__44__29__in1[24]), .B(inst_cellmath__44__29__in0));
INVX2 inst_cellmath__44__29__I1 (.Y(inst_cellmath__44__29__out0[0]), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw3815070899_bdw (
	inst_cellmath__44__28__out0,
	inst_cellmath__44__28__in0,
	inst_cellmath__44__28__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__28__out0;
input [0:0] inst_cellmath__44__28__in0;
input  inst_cellmath__44__28__in1;
wire N5;
NAND2X2 inst_cellmath__44__28__I0 (.Y(N5), .A(inst_cellmath__44__28__in1), .B(inst_cellmath__44__28__in0[0]));
INVX2 inst_cellmath__44__28__I1 (.Y(inst_cellmath__44__28__out0[0]), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw3815070899_bdw (
	inst_cellmath__44__27__out0,
	inst_cellmath__44__27__in0,
	inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__27__out0;
input  inst_cellmath__44__27__in0;
input [0:0] inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3;
wire N7,N8,N9,N10,N11;
NOR2XL inst_cellmath__44__27__I0 (.Y(N7), .A(inst_cellmath__44__27__in0), .B(inst_cellmath__44__27__in2[0]));
INVXL inst_cellmath__44__27__I1 (.Y(N8), .A(N7));
NOR2XL inst_cellmath__44__27__I2 (.Y(N9), .A(N8), .B(inst_cellmath__44__27__in1[0]));
INVXL inst_cellmath__44__27__I3 (.Y(N10), .A(N9));
NOR2X4 inst_cellmath__44__27__I4 (.Y(N11), .A(N10), .B(inst_cellmath__44__27__in3[0]));
INVX2 inst_cellmath__44__27__I5 (.Y(inst_cellmath__44__27__out0[0]), .A(N11));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw3815070899_bdw (
	inst_cellmath__44__26__out0,
	inst_cellmath__44__26__in0,
	inst_cellmath__44__26__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__26__out0;
input [0:0] inst_cellmath__44__26__in0;
input [23:23] inst_cellmath__44__26__in1;
wire N19;
NAND2X4 inst_cellmath__44__26__I4 (.Y(N19), .A(inst_cellmath__44__26__in1[23]), .B(inst_cellmath__44__26__in0[0]));
INVX2 inst_cellmath__44__26__I5 (.Y(inst_cellmath__44__26__out0[0]), .A(N19));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw3815070899_bdw (
	inst_cellmath__44__33__out0,
	inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__33__out0;
input [0:0] inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1;
OR2XL inst_cellmath__44__33__I0 (.Y(inst_cellmath__44__33__out0[0]), .A(inst_cellmath__44__33__in1[0]), .B(inst_cellmath__44__33__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw3815070899_bdw (
	inst_cellmath__44__32__out0,
	inst_cellmath__44__32__in0,
	inst_cellmath__44__32__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__32__out0;
input [0:0] inst_cellmath__44__32__in0;
input  inst_cellmath__44__32__in1;
AND2X1 inst_cellmath__44__32__I0 (.Y(inst_cellmath__44__32__out0[0]), .A(inst_cellmath__44__32__in1), .B(inst_cellmath__44__32__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw3815070899_bdw (
	inst_cellmath__44_0_out0,
	inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__44_0_out0;
input [0:0] inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1;
wire N5;
NOR2X2 inst_cellmath__44_0_I0 (.Y(N5), .A(inst_cellmath__44_0_in0[0]), .B(inst_cellmath__44_0_in1[0]));
INVX2 inst_cellmath__44_0_I1 (.Y(inst_cellmath__44_0_out0), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw3815070899_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__46_0_out0;
input [24:24] inst_cellmath__46_0_in0;
input  inst_cellmath__46_0_in1;
wire N5;
NAND2X2 inst_cellmath__46_0_I0 (.Y(N5), .A(inst_cellmath__46_0_in0[24]), .B(inst_cellmath__46_0_in1));
INVX2 inst_cellmath__46_0_I1 (.Y(inst_cellmath__46_0_out0), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw3815070899_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0;
input [47:47] inst_cellmath__38_0_in1;
wire N5;
NOR2X2 inst_cellmath__38_0_I0 (.Y(N5), .A(inst_cellmath__38_0_in1[47]), .B(inst_cellmath__38_0_in0));
INVX2 inst_cellmath__38_0_I1 (.Y(inst_cellmath__38_0_out0), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw3815070899_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__30_0_out0;
input [7:0] inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
wire N106,N113,N114,N115,N116,N117,N118 
	,N119,N120,N121,N122,N123,N124,N125,N126 
	,N130,N135,N136,N139,N140,N143,N144,N149 
	,N152,N156,N157,N162,N164,N185,N188,N191 
	,N194,N197,N200,N203,N214,N215,N217,N218 
	,N220,N221,N223,N224,N226,N346,N348,N351 
	,N360,N361,N363,N367;
INVXL inst_cellmath__30_0_I40 (.Y(N106), .A(inst_cellmath__30_0_in1[7]));
NOR2X1 inst_cellmath__30_0_I43 (.Y(N113), .A(inst_cellmath__30_0_in1[1]), .B(inst_cellmath__30_0_in0[1]));
NAND2X1 inst_cellmath__30_0_I44 (.Y(N114), .A(inst_cellmath__30_0_in1[1]), .B(inst_cellmath__30_0_in0[1]));
NOR2X1 inst_cellmath__30_0_I45 (.Y(N115), .A(inst_cellmath__30_0_in1[2]), .B(inst_cellmath__30_0_in0[2]));
NAND2X1 inst_cellmath__30_0_I46 (.Y(N116), .A(inst_cellmath__30_0_in1[2]), .B(inst_cellmath__30_0_in0[2]));
NOR2X1 inst_cellmath__30_0_I47 (.Y(N117), .A(inst_cellmath__30_0_in1[3]), .B(inst_cellmath__30_0_in0[3]));
NAND2XL inst_cellmath__30_0_I48 (.Y(N118), .A(inst_cellmath__30_0_in1[3]), .B(inst_cellmath__30_0_in0[3]));
NOR2XL inst_cellmath__30_0_I49 (.Y(N119), .A(inst_cellmath__30_0_in1[4]), .B(inst_cellmath__30_0_in0[4]));
NAND2X1 inst_cellmath__30_0_I50 (.Y(N120), .A(inst_cellmath__30_0_in1[4]), .B(inst_cellmath__30_0_in0[4]));
NOR2XL inst_cellmath__30_0_I51 (.Y(N121), .A(inst_cellmath__30_0_in1[5]), .B(inst_cellmath__30_0_in0[5]));
NAND2XL inst_cellmath__30_0_I52 (.Y(N122), .A(inst_cellmath__30_0_in1[5]), .B(inst_cellmath__30_0_in0[5]));
NOR2XL inst_cellmath__30_0_I53 (.Y(N123), .A(inst_cellmath__30_0_in1[6]), .B(inst_cellmath__30_0_in0[6]));
NAND2XL inst_cellmath__30_0_I54 (.Y(N124), .A(inst_cellmath__30_0_in1[6]), .B(inst_cellmath__30_0_in0[6]));
NOR2XL inst_cellmath__30_0_I55 (.Y(N125), .A(inst_cellmath__30_0_in0[7]), .B(N106));
NAND2XL inst_cellmath__30_0_I56 (.Y(N126), .A(inst_cellmath__30_0_in0[7]), .B(N106));
INVXL inst_cellmath__30_0_I185 (.Y(N346), .A(inst_cellmath__30_0_in1[0]));
INVXL inst_cellmath__30_0_I187 (.Y(N348), .A(inst_cellmath__30_0_in0[0]));
NAND2X2 inst_cellmath__30_0_I60 (.Y(N130), .A(N348), .B(N346));
INVXL inst_cellmath__30_0_I190 (.Y(N351), .A(N113));
AOI21X1 inst_cellmath__30_0_I64 (.Y(N135), .A0(N116), .A1(N113), .B0(N115));
NAND2X1 inst_cellmath__30_0_I65 (.Y(N136), .A(N116), .B(N114));
AOI21XL inst_cellmath__30_0_I68 (.Y(N139), .A0(N120), .A1(N117), .B0(N119));
NAND2XL inst_cellmath__30_0_I69 (.Y(N140), .A(N120), .B(N118));
AOI21XL inst_cellmath__30_0_I72 (.Y(N143), .A0(N124), .A1(N121), .B0(N123));
NAND2XL inst_cellmath__30_0_I73 (.Y(N144), .A(N124), .B(N122));
NAND2XL inst_cellmath__30_0_I76 (.Y(N226), .A(N106), .B(N125));
NAND2XL inst_cellmath__30_0_I77 (.Y(N149), .A(N106), .B(N126));
OAI21X2 inst_cellmath__30_0_I80 (.Y(N152), .A0(N136), .A1(N130), .B0(N135));
INVXL inst_cellmath__30_0_I199 (.Y(N360), .A(N139));
INVXL inst_cellmath__30_0_I200 (.Y(N361), .A(N140));
OAI21XL inst_cellmath__30_0_I84 (.Y(N156), .A0(N144), .A1(N139), .B0(N143));
NOR2XL inst_cellmath__30_0_I85 (.Y(N157), .A(N144), .B(N140));
INVXL inst_cellmath__30_0_I202 (.Y(N363), .A(N152));
AOI21XL inst_cellmath__30_0_I90 (.Y(N162), .A0(N361), .A1(N152), .B0(N360));
AOI21X1 inst_cellmath__30_0_I92 (.Y(N164), .A0(N157), .A1(N152), .B0(N156));
NAND2BXL inst_cellmath__30_0_I112 (.Y(N185), .AN(N113), .B(N114));
NAND2BXL inst_cellmath__30_0_I115 (.Y(N188), .AN(N115), .B(N116));
NAND2BXL inst_cellmath__30_0_I118 (.Y(N191), .AN(N117), .B(N118));
NAND2BXL inst_cellmath__30_0_I121 (.Y(N194), .AN(N119), .B(N120));
NAND2BXL inst_cellmath__30_0_I124 (.Y(N197), .AN(N121), .B(N122));
NAND2BXL inst_cellmath__30_0_I127 (.Y(N200), .AN(N123), .B(N124));
NAND2BXL inst_cellmath__30_0_I130 (.Y(N203), .AN(N125), .B(N126));
INVXL inst_cellmath__30_0_I206 (.Y(N367), .A(N106));
XNOR2X1 inst_cellmath__30_0_I219 (.Y(inst_cellmath__30_0_out0[0]), .A(N346), .B(N348));
XNOR2X1 inst_cellmath__30_0_I209 (.Y(inst_cellmath__30_0_out0[1]), .A(N130), .B(N185));
XNOR2X1 inst_cellmath__30_0_I137 (.Y(inst_cellmath__30_0_out0[3]), .A(N363), .B(N191));
XNOR2X1 inst_cellmath__30_0_I138 (.Y(inst_cellmath__30_0_out0[5]), .A(N162), .B(N197));
XNOR2X1 inst_cellmath__30_0_I139 (.Y(inst_cellmath__30_0_out0[7]), .A(N164), .B(N203));
XOR2XL node_cs_reduced_ii_local_A_I210 (.Y(N215), .A(N188), .B(N114));
XNOR2XL node_cs_reduced_ii_local_A_I167 (.Y(N214), .A(N188), .B(N351));
MX2XL inst_cellmath__30_0_I141 (.Y(inst_cellmath__30_0_out0[2]), .A(N215), .B(N214), .S0(N130));
XOR2XL node_cs_reduced_ii_local_A_I212 (.Y(N218), .A(N194), .B(N118));
XOR2XL node_cs_reduced_ii_local_A_I213 (.Y(N217), .A(N194), .B(N117));
MX2XL inst_cellmath__30_0_I143 (.Y(inst_cellmath__30_0_out0[4]), .A(N218), .B(N217), .S0(N363));
XOR2XL node_cs_reduced_ii_local_A_I214 (.Y(N221), .A(N200), .B(N122));
XOR2XL node_cs_reduced_ii_local_A_I215 (.Y(N220), .A(N200), .B(N121));
MX2XL inst_cellmath__30_0_I145 (.Y(inst_cellmath__30_0_out0[6]), .A(N221), .B(N220), .S0(N162));
XOR2XL node_cs_reduced_ii_local_A_I216 (.Y(N224), .A(N367), .B(N126));
XOR2XL node_cs_reduced_ii_local_A_I217 (.Y(N223), .A(N367), .B(N125));
MX2XL inst_cellmath__30_0_I147 (.Y(inst_cellmath__30_0_out0[8]), .A(N224), .B(N223), .S0(N164));
OAI21XL inst_cellmath__30_0_I225 (.Y(inst_cellmath__30_0_out0[9]), .A0(N149), .A1(N164), .B0(N226));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw3815070899_bdw (
	inst_cellmath__31_0_out0,
	inst_cellmath__31_0_in0
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__31_0_out0;
input [9:0] inst_cellmath__31_0_in0;
wire N77,N116,N121,N127,N132,N135,N141 
	,N197,N201,N294,N439,N443,N446,N450,N467 
	;
INVXL inst_cellmath__31_0_I163 (.Y(inst_cellmath__31_0_out0[0]), .A(inst_cellmath__31_0_in0[0]));
NOR2BX1 inst_cellmath__31_0_I189 (.Y(N77), .AN(inst_cellmath__31_0_in0[1]), .B(inst_cellmath__31_0_out0[0]));
CLKAND2X3 inst_cellmath__31_0_I38 (.Y(N116), .A(inst_cellmath__31_0_in0[2]), .B(N77));
XNOR2X1 inst_cellmath__31_0_I55 (.Y(inst_cellmath__31_0_out0[1]), .A(inst_cellmath__31_0_out0[0]), .B(inst_cellmath__31_0_in0[1]));
XOR2XL inst_cellmath__31_0_I190 (.Y(inst_cellmath__31_0_out0[2]), .A(N77), .B(inst_cellmath__31_0_in0[2]));
NAND2X1 inst_cellmath__31_0_I62 (.Y(N121), .A(inst_cellmath__31_0_in0[3]), .B(N116));
INVXL inst_cellmath__31_0_I173 (.Y(N439), .A(inst_cellmath__31_0_in0[4]));
NAND2X1 inst_cellmath__31_0_I67 (.Y(N127), .A(inst_cellmath__31_0_in0[5]), .B(inst_cellmath__31_0_in0[4]));
NOR2XL inst_cellmath__31_0_I72 (.Y(N132), .A(N439), .B(N121));
NOR2X2 inst_cellmath__31_0_I74 (.Y(N135), .A(N127), .B(N121));
INVXL inst_cellmath__31_0_I177 (.Y(N443), .A(inst_cellmath__31_0_in0[6]));
NAND2X1 inst_cellmath__31_0_I79 (.Y(N141), .A(inst_cellmath__31_0_in0[7]), .B(inst_cellmath__31_0_in0[6]));
INVXL inst_cellmath__31_0_I180 (.Y(N446), .A(inst_cellmath__31_0_in0[8]));
NOR2XL inst_cellmath__31_0_I89 (.Y(N294), .A(N446), .B(N141));
INVXL inst_cellmath__31_0_I184 (.Y(N450), .A(inst_cellmath__31_0_in0[7]));
XOR2XL inst_cellmath__31_0_I193 (.Y(inst_cellmath__31_0_out0[3]), .A(N116), .B(inst_cellmath__31_0_in0[3]));
XOR2XL inst_cellmath__31_0_I282 (.Y(inst_cellmath__31_0_out0[4]), .A(N121), .B(N439));
XOR2XL inst_cellmath__31_0_I277 (.Y(inst_cellmath__31_0_out0[5]), .A(N132), .B(inst_cellmath__31_0_in0[5]));
XNOR2XL inst_cellmath__31_0_I278 (.Y(inst_cellmath__31_0_out0[6]), .A(N135), .B(N443));
XNOR2XL inst_cellmath__31_0_I279 (.Y(N197), .A(N450), .B(N443));
MXI2XL inst_cellmath__31_0_I122 (.Y(inst_cellmath__31_0_out0[7]), .A(N450), .B(N197), .S0(N135));
XNOR2X1 inst_cellmath__31_0_I149 (.Y(N201), .A(N446), .B(N141));
MXI2XL inst_cellmath__31_0_I124 (.Y(inst_cellmath__31_0_out0[8]), .A(N446), .B(N201), .S0(N135));
NAND2XL node_cs_const1_cs_ii_A_I210 (.Y(N467), .A(N294), .B(N135));
XNOR2X1 node_cs_const1_cs_ii_A_I280 (.Y(inst_cellmath__31_0_out0[9]), .A(inst_cellmath__31_0_in0[9]), .B(N467));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw3815070899_bdw (
	inst_cellmath__48_0_out0,
	inst_cellmath__48_0_in0,
	inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__48_0_out0;
input  inst_cellmath__48_0_in0;
input [9:0] inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2;
wire N33,N34,N35,N36,N37,N38,N39 
	,N40,N41,N42,N43,N44,N45,N46,N47 
	,N48,N49,N50,N51,N52;
INVXL inst_cellmath__48_0_I0 (.Y(N33), .A(inst_cellmath__48_0_in1[0]));
INVXL inst_cellmath__48_0_I1 (.Y(N34), .A(inst_cellmath__48_0_in1[1]));
INVXL inst_cellmath__48_0_I2 (.Y(N35), .A(inst_cellmath__48_0_in1[2]));
INVXL inst_cellmath__48_0_I3 (.Y(N36), .A(inst_cellmath__48_0_in1[3]));
INVXL inst_cellmath__48_0_I4 (.Y(N37), .A(inst_cellmath__48_0_in1[4]));
INVXL inst_cellmath__48_0_I5 (.Y(N38), .A(inst_cellmath__48_0_in1[5]));
INVXL inst_cellmath__48_0_I6 (.Y(N39), .A(inst_cellmath__48_0_in1[6]));
INVXL inst_cellmath__48_0_I7 (.Y(N40), .A(inst_cellmath__48_0_in1[7]));
INVXL inst_cellmath__48_0_I8 (.Y(N41), .A(inst_cellmath__48_0_in1[8]));
INVXL inst_cellmath__48_0_I9 (.Y(N42), .A(inst_cellmath__48_0_in1[9]));
INVXL inst_cellmath__48_0_I10 (.Y(N43), .A(inst_cellmath__48_0_in2[0]));
INVXL inst_cellmath__48_0_I11 (.Y(N44), .A(inst_cellmath__48_0_in2[1]));
INVXL inst_cellmath__48_0_I12 (.Y(N45), .A(inst_cellmath__48_0_in2[2]));
INVXL inst_cellmath__48_0_I13 (.Y(N46), .A(inst_cellmath__48_0_in2[3]));
INVXL inst_cellmath__48_0_I14 (.Y(N47), .A(inst_cellmath__48_0_in2[4]));
INVXL inst_cellmath__48_0_I15 (.Y(N48), .A(inst_cellmath__48_0_in2[5]));
INVXL inst_cellmath__48_0_I16 (.Y(N49), .A(inst_cellmath__48_0_in2[6]));
INVXL inst_cellmath__48_0_I17 (.Y(N50), .A(inst_cellmath__48_0_in2[7]));
INVXL inst_cellmath__48_0_I18 (.Y(N51), .A(inst_cellmath__48_0_in2[8]));
INVXL inst_cellmath__48_0_I19 (.Y(N52), .A(inst_cellmath__48_0_in2[9]));
MXI2X1 inst_cellmath__48_0_I20 (.Y(inst_cellmath__48_0_out0[0]), .A(N43), .B(N33), .S0(inst_cellmath__48_0_in0));
MXI2X1 inst_cellmath__48_0_I21 (.Y(inst_cellmath__48_0_out0[1]), .A(N44), .B(N34), .S0(inst_cellmath__48_0_in0));
MXI2XL inst_cellmath__48_0_I22 (.Y(inst_cellmath__48_0_out0[2]), .A(N45), .B(N35), .S0(inst_cellmath__48_0_in0));
MXI2X2 inst_cellmath__48_0_I23 (.Y(inst_cellmath__48_0_out0[3]), .A(N46), .B(N36), .S0(inst_cellmath__48_0_in0));
MXI2X2 inst_cellmath__48_0_I24 (.Y(inst_cellmath__48_0_out0[4]), .A(N47), .B(N37), .S0(inst_cellmath__48_0_in0));
MXI2X2 inst_cellmath__48_0_I25 (.Y(inst_cellmath__48_0_out0[5]), .A(N48), .B(N38), .S0(inst_cellmath__48_0_in0));
MXI2X2 inst_cellmath__48_0_I26 (.Y(inst_cellmath__48_0_out0[6]), .A(N49), .B(N39), .S0(inst_cellmath__48_0_in0));
MXI2X2 inst_cellmath__48_0_I27 (.Y(inst_cellmath__48_0_out0[7]), .A(N50), .B(N40), .S0(inst_cellmath__48_0_in0));
MXI2XL inst_cellmath__48_0_I28 (.Y(inst_cellmath__48_0_out0[8]), .A(N51), .B(N41), .S0(inst_cellmath__48_0_in0));
MXI2XL inst_cellmath__48_0_I29 (.Y(inst_cellmath__48_0_out0[9]), .A(N52), .B(N42), .S0(inst_cellmath__48_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw3815070899_bdw (
	inst_cellmath__51__49__out0,
	inst_cellmath__51__49__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__49__out0;
input [7:0] inst_cellmath__51__49__in0;
wire N11,N12,N13,N14,N15,N16,N17 
	;
NAND2X2 inst_cellmath__51__49__I0 (.Y(N11), .A(inst_cellmath__51__49__in0[0]), .B(inst_cellmath__51__49__in0[1]));
NAND2X4 inst_cellmath__51__49__I1 (.Y(N12), .A(inst_cellmath__51__49__in0[7]), .B(inst_cellmath__51__49__in0[6]));
NAND2X4 inst_cellmath__51__49__I2 (.Y(N13), .A(inst_cellmath__51__49__in0[5]), .B(inst_cellmath__51__49__in0[4]));
NAND2X4 inst_cellmath__51__49__I3 (.Y(N14), .A(inst_cellmath__51__49__in0[3]), .B(inst_cellmath__51__49__in0[2]));
NOR2X4 inst_cellmath__51__49__I4 (.Y(N15), .A(N11), .B(N12));
NOR2X4 inst_cellmath__51__49__I5 (.Y(N16), .A(N13), .B(N14));
NAND2X2 inst_cellmath__51__49__I6 (.Y(N17), .A(N15), .B(N16));
INVX1 inst_cellmath__51__49__I7 (.Y(inst_cellmath__51__49__out0[0]), .A(N17));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw3815070899_bdw (
	inst_cellmath__51__48__out0,
	inst_cellmath__51__48__in0,
	inst_cellmath__51__48__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__48__out0;
input [0:0] inst_cellmath__51__48__in0;
input [8:8] inst_cellmath__51__48__in1;
wire N5;
NOR2X2 inst_cellmath__51__48__I0 (.Y(N5), .A(inst_cellmath__51__48__in1[8]), .B(inst_cellmath__51__48__in0[0]));
INVX2 inst_cellmath__51__48__I1 (.Y(inst_cellmath__51__48__out0[0]), .A(N5));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw3815070899_bdw (
	inst_cellmath__51_0_out0,
	inst_cellmath__51_0_in0,
	inst_cellmath__51_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__51_0_out0;
input [0:0] inst_cellmath__51_0_in0;
input [9:9] inst_cellmath__51_0_in1;
wire N5;
INVXL inst_cellmath__51_0_I0 (.Y(N5), .A(inst_cellmath__51_0_in1[9]));
CLKAND2X6 inst_cellmath__51_0_I1 (.Y(inst_cellmath__51_0_out0), .A(N5), .B(inst_cellmath__51_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw3815070899_bdw (
	inst_cellmath__28_0_out0,
	inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__28_0_out0;
input  inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1;
wire N19;
NOR2X2 inst_cellmath__28_0_I4 (.Y(N19), .A(inst_cellmath__28_0_in0), .B(inst_cellmath__28_0_in1));
INVX1 inst_cellmath__28_0_I5 (.Y(inst_cellmath__28_0_out0), .A(N19));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw3815070899_bdw (
	inst_cellmath__27_0_out0,
	inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__27_0_out0;
input  inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1;
OR2XL inst_cellmath__27_0_I0 (.Y(inst_cellmath__27_0_out0), .A(inst_cellmath__27_0_in0), .B(inst_cellmath__27_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw3815070899_bdw (
	inst_cellmath__50__50__out0,
	inst_cellmath__50__50__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__50__50__out0;
input [9:0] inst_cellmath__50__50__in0;
wire N13,N14,N15,N16,N18,N20,N21 
	,N22;
NOR2XL inst_cellmath__50__50__I0 (.Y(N13), .A(inst_cellmath__50__50__in0[9]), .B(inst_cellmath__50__50__in0[1]));
NOR2X1 inst_cellmath__50__50__I1 (.Y(N14), .A(inst_cellmath__50__50__in0[2]), .B(inst_cellmath__50__50__in0[6]));
NOR2X1 inst_cellmath__50__50__I2 (.Y(N15), .A(inst_cellmath__50__50__in0[4]), .B(inst_cellmath__50__50__in0[8]));
NOR2X4 inst_cellmath__50__50__I3 (.Y(N16), .A(inst_cellmath__50__50__in0[7]), .B(inst_cellmath__50__50__in0[5]));
NAND2X1 inst_cellmath__50__50__I5 (.Y(N18), .A(N13), .B(N14));
OR2XL inst_cellmath__50__50__I77 (.Y(N20), .A(inst_cellmath__50__50__in0[3]), .B(inst_cellmath__50__50__in0[0]));
NOR2X1 inst_cellmath__50__50__I8 (.Y(N21), .A(N20), .B(N18));
CLKAND2X2 inst_cellmath__50__50__I79 (.Y(N22), .A(N15), .B(N16));
NAND2X2 inst_cellmath__50__50__I10 (.Y(inst_cellmath__50__50__out0[0]), .A(N22), .B(N21));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw3815070899_bdw (
	inst_cellmath__49_1_out0,
	inst_cellmath__49_1_in0,
	inst_cellmath__49_1_in1,
	inst_cellmath__49_1_in2,
	inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__49_1_out0;
input  inst_cellmath__49_1_in0;
input [0:0] inst_cellmath__49_1_in1;
input [9:9] inst_cellmath__49_1_in2;
input  inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5;
wire N9,N10,N11,N12,N13,N14,N15 
	;
NOR2XL inst_cellmath__49_1_I0 (.Y(N9), .A(inst_cellmath__49_1_in3), .B(inst_cellmath__49_1_in4));
INVXL inst_cellmath__49_1_I1 (.Y(N10), .A(N9));
NOR2XL inst_cellmath__49_1_I2 (.Y(N11), .A(N10), .B(inst_cellmath__49_1_in5));
INVXL inst_cellmath__49_1_I3 (.Y(N12), .A(N11));
NOR2XL inst_cellmath__49_1_I4 (.Y(N13), .A(N12), .B(inst_cellmath__49_1_in2[9]));
NAND2X2 inst_cellmath__49_1_I5 (.Y(N14), .A(N13), .B(inst_cellmath__49_1_in1[0]));
NOR2X4 inst_cellmath__49_1_I6 (.Y(N15), .A(N14), .B(inst_cellmath__49_1_in0));
CLKINVX4 inst_cellmath__49_1_I7 (.Y(inst_cellmath__49_1_out0), .A(N15));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw3815070899_bdw (
	inst_cellmath__37__43__out0,
	inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__43__out0;
input  inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1;
OR2XL inst_cellmath__37__43__I0 (.Y(inst_cellmath__37__43__out0[0]), .A(inst_cellmath__37__43__in0), .B(inst_cellmath__37__43__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw3815070899_bdw (
	inst_cellmath__32__11__out0,
	inst_cellmath__32__11__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__32__11__out0;
input [8:7] inst_cellmath__32__11__in0;
wire N21;
NOR2XL inst_cellmath__32__11__I5 (.Y(N21), .A(inst_cellmath__32__11__in0[8]), .B(inst_cellmath__32__11__in0[7]));
INVXL inst_cellmath__32__11__I6 (.Y(inst_cellmath__32__11__out0[0]), .A(N21));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw3815070899_bdw (
	inst_cellmath__32__10__out0,
	inst_cellmath__32__10__in0,
	inst_cellmath__32__10__in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__32__10__out0;
input [0:0] inst_cellmath__32__10__in0;
input [9:9] inst_cellmath__32__10__in1;
wire N5;
INVXL inst_cellmath__32__10__I0 (.Y(N5), .A(inst_cellmath__32__10__in1[9]));
NAND2X2 inst_cellmath__32__10__I1 (.Y(inst_cellmath__32__10__out0), .A(N5), .B(inst_cellmath__32__10__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw3815070899_bdw (
	inst_cellmath__37__42__out0,
	inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__42__out0;
input  inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1;
OR2XL inst_cellmath__37__42__I0 (.Y(inst_cellmath__37__42__out0[0]), .A(inst_cellmath__37__42__in1), .B(inst_cellmath__37__42__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw3815070899_bdw (
	inst_cellmath__7_0_out0,
	inst_cellmath__7_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__7_0_out0;
input [2:0] inst_cellmath__7_0_in0;
wire N36,N38;
INVX1 inst_cellmath__7_0_I19 (.Y(N36), .A(inst_cellmath__7_0_in0[2]));
NAND3X1 inst_cellmath__7_0_I20 (.Y(N38), .A(inst_cellmath__7_0_in0[0]), .B(inst_cellmath__7_0_in0[1]), .C(N36));
INVXL inst_cellmath__7_0_I21 (.Y(inst_cellmath__7_0_out0), .A(N38));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw3815070899_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__42_0_out0;
input  inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3;
wire N9,N12;
INVXL inst_cellmath__42_0_I0 (.Y(N9), .A(inst_cellmath__42_0_in0));
MXI2XL inst_cellmath__42_0_I3 (.Y(N12), .A(N9), .B(inst_cellmath__42_0_in3), .S0(inst_cellmath__42_0_in1));
MXI2XL inst_cellmath__42_0_I4 (.Y(inst_cellmath__42_0_out0), .A(N12), .B(inst_cellmath__42_0_in3), .S0(inst_cellmath__42_0_in2));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw3815070899_bdw (
	inst_cellmath__52_0_out0,
	inst_cellmath__52_0_in0,
	inst_cellmath__52_0_in1,
	inst_cellmath__52_0_in2,
	inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__52_0_out0;
input  inst_cellmath__52_0_in0;
input [7:0] inst_cellmath__52_0_in1;
input  inst_cellmath__52_0_in2;
input [0:0] inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4;
wire N41,N50,N66,N67,N68,N69,N70 
	,N71,N72,N73,N82;
NOR2BX1 inst_cellmath__52_0_I197 (.Y(N41), .AN(inst_cellmath__52_0_in2), .B(inst_cellmath__52_0_in4[0]));
NOR2XL inst_cellmath__52_0_I16 (.Y(N50), .A(N41), .B(inst_cellmath__52_0_in3[0]));
NOR2BX1 inst_cellmath__52_0_I198 (.Y(N82), .AN(inst_cellmath__52_0_in4[0]), .B(inst_cellmath__52_0_in3[0]));
INVXL inst_cellmath__52_0_I24 (.Y(N66), .A(inst_cellmath__52_0_in1[0]));
INVXL inst_cellmath__52_0_I25 (.Y(N67), .A(inst_cellmath__52_0_in1[1]));
INVXL inst_cellmath__52_0_I26 (.Y(N68), .A(inst_cellmath__52_0_in1[2]));
INVXL inst_cellmath__52_0_I27 (.Y(N69), .A(inst_cellmath__52_0_in1[3]));
INVXL inst_cellmath__52_0_I28 (.Y(N70), .A(inst_cellmath__52_0_in1[4]));
INVXL inst_cellmath__52_0_I29 (.Y(N71), .A(inst_cellmath__52_0_in1[5]));
INVXL inst_cellmath__52_0_I30 (.Y(N72), .A(inst_cellmath__52_0_in1[6]));
INVXL inst_cellmath__52_0_I31 (.Y(N73), .A(inst_cellmath__52_0_in1[7]));
MXI2XL inst_cellmath__52_0_I32 (.Y(inst_cellmath__52_0_out0[0]), .A(N66), .B(N50), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I33 (.Y(inst_cellmath__52_0_out0[1]), .A(N67), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I34 (.Y(inst_cellmath__52_0_out0[2]), .A(N68), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I35 (.Y(inst_cellmath__52_0_out0[3]), .A(N69), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I36 (.Y(inst_cellmath__52_0_out0[4]), .A(N70), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I37 (.Y(inst_cellmath__52_0_out0[5]), .A(N71), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I38 (.Y(inst_cellmath__52_0_out0[6]), .A(N72), .B(N82), .S0(inst_cellmath__52_0_in0));
MXI2XL inst_cellmath__52_0_I39 (.Y(inst_cellmath__52_0_out0[7]), .A(N73), .B(N82), .S0(inst_cellmath__52_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw3815070899_bdw (
	inst_cellmath__47_0_out0,
	inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__47_0_out0;
input  inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4;
wire N10,N12;
OR3XL inst_cellmath__47_0_I7 (.Y(N10), .A(inst_cellmath__47_0_in2), .B(inst_cellmath__47_0_in3), .C(inst_cellmath__47_0_in4));
OR2XL inst_cellmath__47_0_I4 (.Y(N12), .A(inst_cellmath__47_0_in0), .B(N10));
NOR2X2 inst_cellmath__47_0_I5 (.Y(inst_cellmath__47_0_out0), .A(N12), .B(inst_cellmath__47_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw3815070899_bdw (
	inst_cellmath__53_U_out0,
	inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1,
	inst_cellmath__53_U_in2,
	inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4,
	inst_cellmath__53_U_in5
	); /* architecture "gate_level" */ 
output [22:22] inst_cellmath__53_U_out0;
input  inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1;
input [22:22] inst_cellmath__53_U_in2;
input  inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4;
input [46:46] inst_cellmath__53_U_in5;
wire N12,N14;
NOR2XL inst_cellmath__53_U_I0 (.Y(N12), .A(inst_cellmath__53_U_in1), .B(inst_cellmath__53_U_in4));
MXI2XL inst_cellmath__53_U_I1 (.Y(N14), .A(inst_cellmath__53_U_in5[46]), .B(inst_cellmath__53_U_in2[22]), .S0(inst_cellmath__53_U_in3));
MXI2XL inst_cellmath__53_U_I2 (.Y(inst_cellmath__53_U_out0[22]), .A(N14), .B(N12), .S0(inst_cellmath__53_U_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw3815070899_bdw (
	inst_cellmath__53_M_out0,
	inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1,
	inst_cellmath__53_M_in2,
	inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4,
	inst_cellmath__53_M_in5,
	inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7,
	inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9
	); /* architecture "gate_level" */ 
output [21:0] inst_cellmath__53_M_out0;
input  inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1;
input [21:0] inst_cellmath__53_M_in2;
input  inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4;
input [45:24] inst_cellmath__53_M_in5;
input  inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7;
input [21:0] inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9;
wire N145,N147,N149,N151,N153,N155,N157 
	,N159,N161,N163,N165,N167,N169,N171,N173 
	,N175,N177,N179,N181,N183,N185,N187,N189 
	,N190,N191,N192,N193,N194,N195,N196,N197 
	,N198,N199,N200,N201,N202,N203,N204,N205 
	,N206,N207,N208,N209,N210,N211,N212,N213 
	,N214,N215,N216,N217,N218,N219,N220,N221 
	,N222,N223,N224,N225,N226,N227,N228,N229 
	,N230,N231,N232,N233,N234,N235,N236,N237 
	,N238,N239,N240,N241,N242,N243,N244,N245 
	,N246,N247,N248,N249,N250,N251,N252,N253 
	,N254,N377,N378,N384,N390,N396,N398,N404 
	,N407,N412,N417,N422,N427;
INVXL buf1_A_I181 (.Y(N422), .A(inst_cellmath__53_M_in6));
INVXL buf1_A_I182 (.Y(N398), .A(N422));
AND2XL inst_cellmath__53_M_I22 (.Y(N145), .A(inst_cellmath__53_M_in8[0]), .B(N398));
AND2XL inst_cellmath__53_M_I23 (.Y(N147), .A(inst_cellmath__53_M_in8[1]), .B(N398));
AND2XL inst_cellmath__53_M_I24 (.Y(N149), .A(inst_cellmath__53_M_in8[2]), .B(N398));
AND2XL inst_cellmath__53_M_I25 (.Y(N151), .A(inst_cellmath__53_M_in8[3]), .B(N398));
AND2XL inst_cellmath__53_M_I26 (.Y(N153), .A(inst_cellmath__53_M_in8[4]), .B(N398));
AND2XL inst_cellmath__53_M_I27 (.Y(N155), .A(inst_cellmath__53_M_in8[5]), .B(N398));
AND2XL inst_cellmath__53_M_I28 (.Y(N157), .A(inst_cellmath__53_M_in8[6]), .B(N398));
AND2XL inst_cellmath__53_M_I29 (.Y(N159), .A(inst_cellmath__53_M_in8[7]), .B(N398));
AND2XL inst_cellmath__53_M_I30 (.Y(N161), .A(inst_cellmath__53_M_in8[8]), .B(N398));
AND2XL inst_cellmath__53_M_I31 (.Y(N163), .A(inst_cellmath__53_M_in8[9]), .B(N398));
AND2XL inst_cellmath__53_M_I32 (.Y(N165), .A(inst_cellmath__53_M_in8[10]), .B(N398));
AND2XL inst_cellmath__53_M_I33 (.Y(N167), .A(inst_cellmath__53_M_in8[11]), .B(N398));
AND2XL inst_cellmath__53_M_I34 (.Y(N169), .A(inst_cellmath__53_M_in8[12]), .B(N398));
AND2XL inst_cellmath__53_M_I35 (.Y(N171), .A(inst_cellmath__53_M_in8[13]), .B(N398));
AND2XL inst_cellmath__53_M_I36 (.Y(N173), .A(inst_cellmath__53_M_in8[14]), .B(N398));
AND2XL inst_cellmath__53_M_I37 (.Y(N175), .A(inst_cellmath__53_M_in8[15]), .B(N398));
AND2XL inst_cellmath__53_M_I38 (.Y(N177), .A(inst_cellmath__53_M_in8[16]), .B(N398));
AND2XL inst_cellmath__53_M_I39 (.Y(N179), .A(inst_cellmath__53_M_in8[17]), .B(N398));
AND2XL inst_cellmath__53_M_I40 (.Y(N181), .A(inst_cellmath__53_M_in8[18]), .B(N398));
AND2XL inst_cellmath__53_M_I41 (.Y(N183), .A(inst_cellmath__53_M_in8[19]), .B(N398));
AND2XL inst_cellmath__53_M_I42 (.Y(N185), .A(inst_cellmath__53_M_in8[20]), .B(N398));
AND2XL inst_cellmath__53_M_I43 (.Y(N187), .A(inst_cellmath__53_M_in8[21]), .B(N398));
INVXL buf1_A_I183 (.Y(N427), .A(inst_cellmath__53_M_in7));
INVXL buf1_A_I184 (.Y(N404), .A(N427));
MX2XL inst_cellmath__53_M_I44 (.Y(N189), .A(N145), .B(inst_cellmath__53_M_in9[0]), .S0(N404));
MX2XL inst_cellmath__53_M_I45 (.Y(N190), .A(N147), .B(inst_cellmath__53_M_in9[1]), .S0(N404));
MX2XL inst_cellmath__53_M_I46 (.Y(N191), .A(N149), .B(inst_cellmath__53_M_in9[2]), .S0(N404));
MX2XL inst_cellmath__53_M_I47 (.Y(N192), .A(N151), .B(inst_cellmath__53_M_in9[3]), .S0(N404));
MX2XL inst_cellmath__53_M_I48 (.Y(N193), .A(N153), .B(inst_cellmath__53_M_in9[4]), .S0(N404));
MX2XL inst_cellmath__53_M_I49 (.Y(N194), .A(N155), .B(inst_cellmath__53_M_in9[5]), .S0(N404));
MX2XL inst_cellmath__53_M_I50 (.Y(N195), .A(N157), .B(inst_cellmath__53_M_in9[6]), .S0(N404));
MX2XL inst_cellmath__53_M_I51 (.Y(N196), .A(N159), .B(inst_cellmath__53_M_in9[7]), .S0(N404));
MX2XL inst_cellmath__53_M_I52 (.Y(N197), .A(N161), .B(inst_cellmath__53_M_in9[8]), .S0(N404));
MX2XL inst_cellmath__53_M_I53 (.Y(N198), .A(N163), .B(inst_cellmath__53_M_in9[9]), .S0(N404));
MX2XL inst_cellmath__53_M_I54 (.Y(N199), .A(N165), .B(inst_cellmath__53_M_in9[10]), .S0(N404));
MX2XL inst_cellmath__53_M_I55 (.Y(N200), .A(N167), .B(inst_cellmath__53_M_in9[11]), .S0(N404));
MX2XL inst_cellmath__53_M_I56 (.Y(N201), .A(N169), .B(inst_cellmath__53_M_in9[12]), .S0(N404));
MX2XL inst_cellmath__53_M_I57 (.Y(N202), .A(N171), .B(inst_cellmath__53_M_in9[13]), .S0(N404));
MX2XL inst_cellmath__53_M_I58 (.Y(N203), .A(N173), .B(inst_cellmath__53_M_in9[14]), .S0(N404));
MX2XL inst_cellmath__53_M_I59 (.Y(N204), .A(N175), .B(inst_cellmath__53_M_in9[15]), .S0(N404));
MX2XL inst_cellmath__53_M_I60 (.Y(N205), .A(N177), .B(inst_cellmath__53_M_in9[16]), .S0(N404));
MX2XL inst_cellmath__53_M_I61 (.Y(N206), .A(N179), .B(inst_cellmath__53_M_in9[17]), .S0(N404));
MX2XL inst_cellmath__53_M_I62 (.Y(N207), .A(N181), .B(inst_cellmath__53_M_in9[18]), .S0(N404));
MX2XL inst_cellmath__53_M_I63 (.Y(N208), .A(N183), .B(inst_cellmath__53_M_in9[19]), .S0(N404));
MX2XL inst_cellmath__53_M_I64 (.Y(N209), .A(N185), .B(inst_cellmath__53_M_in9[20]), .S0(N404));
MX2XL inst_cellmath__53_M_I65 (.Y(N210), .A(N187), .B(inst_cellmath__53_M_in9[21]), .S0(N404));
INVXL buf1_A_I175 (.Y(N407), .A(inst_cellmath__53_M_in1));
INVXL buf1_A_I176 (.Y(N384), .A(N407));
INVXL buf1_A_I179 (.Y(N417), .A(inst_cellmath__53_M_in4));
INVXL buf1_A_I180 (.Y(N396), .A(N417));
MXI2XL inst_cellmath__53_M_I66 (.Y(N211), .A(N384), .B(N189), .S0(N396));
MXI2XL inst_cellmath__53_M_I67 (.Y(N212), .A(N384), .B(N190), .S0(N396));
MXI2XL inst_cellmath__53_M_I68 (.Y(N213), .A(N384), .B(N191), .S0(N396));
MXI2XL inst_cellmath__53_M_I69 (.Y(N214), .A(N384), .B(N192), .S0(N396));
MXI2XL inst_cellmath__53_M_I70 (.Y(N215), .A(N384), .B(N193), .S0(N396));
MXI2XL inst_cellmath__53_M_I71 (.Y(N216), .A(N384), .B(N194), .S0(N396));
MXI2XL inst_cellmath__53_M_I72 (.Y(N217), .A(N384), .B(N195), .S0(N396));
MXI2XL inst_cellmath__53_M_I73 (.Y(N218), .A(N384), .B(N196), .S0(N396));
MXI2XL inst_cellmath__53_M_I74 (.Y(N219), .A(N384), .B(N197), .S0(N396));
MXI2XL inst_cellmath__53_M_I75 (.Y(N220), .A(N384), .B(N198), .S0(N396));
MXI2XL inst_cellmath__53_M_I76 (.Y(N221), .A(N384), .B(N199), .S0(N396));
MXI2XL inst_cellmath__53_M_I77 (.Y(N222), .A(N384), .B(N200), .S0(N396));
MXI2XL inst_cellmath__53_M_I78 (.Y(N223), .A(N384), .B(N201), .S0(N396));
MXI2XL inst_cellmath__53_M_I79 (.Y(N224), .A(N384), .B(N202), .S0(N396));
MXI2XL inst_cellmath__53_M_I80 (.Y(N225), .A(N384), .B(N203), .S0(N396));
MXI2XL inst_cellmath__53_M_I81 (.Y(N226), .A(N384), .B(N204), .S0(N396));
MXI2XL inst_cellmath__53_M_I82 (.Y(N227), .A(N384), .B(N205), .S0(N396));
MXI2XL inst_cellmath__53_M_I83 (.Y(N228), .A(N384), .B(N206), .S0(N396));
MXI2XL inst_cellmath__53_M_I84 (.Y(N229), .A(N384), .B(N207), .S0(N396));
MXI2XL inst_cellmath__53_M_I85 (.Y(N230), .A(N384), .B(N208), .S0(N396));
MXI2XL inst_cellmath__53_M_I86 (.Y(N231), .A(N384), .B(N209), .S0(N396));
MXI2XL inst_cellmath__53_M_I87 (.Y(N232), .A(N384), .B(N210), .S0(N396));
INVXL buf1_A_I177 (.Y(N412), .A(inst_cellmath__53_M_in3));
INVXL buf1_A_I178 (.Y(N390), .A(N412));
MXI2XL inst_cellmath__53_M_I88 (.Y(N233), .A(inst_cellmath__53_M_in5[24]), .B(inst_cellmath__53_M_in2[0]), .S0(N390));
MXI2XL inst_cellmath__53_M_I89 (.Y(N234), .A(inst_cellmath__53_M_in5[25]), .B(inst_cellmath__53_M_in2[1]), .S0(N390));
MXI2XL inst_cellmath__53_M_I90 (.Y(N235), .A(inst_cellmath__53_M_in5[26]), .B(inst_cellmath__53_M_in2[2]), .S0(N390));
MXI2XL inst_cellmath__53_M_I91 (.Y(N236), .A(inst_cellmath__53_M_in5[27]), .B(inst_cellmath__53_M_in2[3]), .S0(N390));
MXI2XL inst_cellmath__53_M_I92 (.Y(N237), .A(inst_cellmath__53_M_in5[28]), .B(inst_cellmath__53_M_in2[4]), .S0(N390));
MXI2XL inst_cellmath__53_M_I93 (.Y(N238), .A(inst_cellmath__53_M_in5[29]), .B(inst_cellmath__53_M_in2[5]), .S0(N390));
MXI2XL inst_cellmath__53_M_I94 (.Y(N239), .A(inst_cellmath__53_M_in5[30]), .B(inst_cellmath__53_M_in2[6]), .S0(N390));
MXI2XL inst_cellmath__53_M_I95 (.Y(N240), .A(inst_cellmath__53_M_in5[31]), .B(inst_cellmath__53_M_in2[7]), .S0(N390));
MXI2XL inst_cellmath__53_M_I96 (.Y(N241), .A(inst_cellmath__53_M_in5[32]), .B(inst_cellmath__53_M_in2[8]), .S0(N390));
MXI2XL inst_cellmath__53_M_I97 (.Y(N242), .A(inst_cellmath__53_M_in5[33]), .B(inst_cellmath__53_M_in2[9]), .S0(N390));
MXI2XL inst_cellmath__53_M_I98 (.Y(N243), .A(inst_cellmath__53_M_in5[34]), .B(inst_cellmath__53_M_in2[10]), .S0(N390));
MXI2XL inst_cellmath__53_M_I99 (.Y(N244), .A(inst_cellmath__53_M_in5[35]), .B(inst_cellmath__53_M_in2[11]), .S0(N390));
MXI2XL inst_cellmath__53_M_I100 (.Y(N245), .A(inst_cellmath__53_M_in5[36]), .B(inst_cellmath__53_M_in2[12]), .S0(N390));
MXI2XL inst_cellmath__53_M_I101 (.Y(N246), .A(inst_cellmath__53_M_in5[37]), .B(inst_cellmath__53_M_in2[13]), .S0(N390));
MXI2XL inst_cellmath__53_M_I102 (.Y(N247), .A(inst_cellmath__53_M_in5[38]), .B(inst_cellmath__53_M_in2[14]), .S0(N390));
MXI2XL inst_cellmath__53_M_I103 (.Y(N248), .A(inst_cellmath__53_M_in5[39]), .B(inst_cellmath__53_M_in2[15]), .S0(N390));
MXI2XL inst_cellmath__53_M_I104 (.Y(N249), .A(inst_cellmath__53_M_in5[40]), .B(inst_cellmath__53_M_in2[16]), .S0(N390));
MXI2XL inst_cellmath__53_M_I105 (.Y(N250), .A(inst_cellmath__53_M_in5[41]), .B(inst_cellmath__53_M_in2[17]), .S0(N390));
MXI2XL inst_cellmath__53_M_I106 (.Y(N251), .A(inst_cellmath__53_M_in5[42]), .B(inst_cellmath__53_M_in2[18]), .S0(N390));
MXI2XL inst_cellmath__53_M_I107 (.Y(N252), .A(inst_cellmath__53_M_in5[43]), .B(inst_cellmath__53_M_in2[19]), .S0(N390));
MXI2XL inst_cellmath__53_M_I108 (.Y(N253), .A(inst_cellmath__53_M_in5[44]), .B(inst_cellmath__53_M_in2[20]), .S0(N390));
MXI2XL inst_cellmath__53_M_I109 (.Y(N254), .A(inst_cellmath__53_M_in5[45]), .B(inst_cellmath__53_M_in2[21]), .S0(N390));
CLKINVX8 inst_cellmath__53_M_I138 (.Y(N377), .A(inst_cellmath__53_M_in0));
CLKINVX8 inst_cellmath__53_M_I139 (.Y(N378), .A(N377));
MXI2XL inst_cellmath__53_M_I110 (.Y(inst_cellmath__53_M_out0[0]), .A(N233), .B(N211), .S0(N378));
MXI2XL inst_cellmath__53_M_I111 (.Y(inst_cellmath__53_M_out0[1]), .A(N234), .B(N212), .S0(N378));
MXI2XL inst_cellmath__53_M_I112 (.Y(inst_cellmath__53_M_out0[2]), .A(N235), .B(N213), .S0(N378));
MXI2XL inst_cellmath__53_M_I113 (.Y(inst_cellmath__53_M_out0[3]), .A(N236), .B(N214), .S0(N378));
MXI2XL inst_cellmath__53_M_I114 (.Y(inst_cellmath__53_M_out0[4]), .A(N237), .B(N215), .S0(N378));
MXI2XL inst_cellmath__53_M_I115 (.Y(inst_cellmath__53_M_out0[5]), .A(N238), .B(N216), .S0(N378));
MXI2XL inst_cellmath__53_M_I116 (.Y(inst_cellmath__53_M_out0[6]), .A(N239), .B(N217), .S0(N378));
MXI2XL inst_cellmath__53_M_I117 (.Y(inst_cellmath__53_M_out0[7]), .A(N240), .B(N218), .S0(N378));
MXI2XL inst_cellmath__53_M_I118 (.Y(inst_cellmath__53_M_out0[8]), .A(N241), .B(N219), .S0(N378));
MXI2XL inst_cellmath__53_M_I119 (.Y(inst_cellmath__53_M_out0[9]), .A(N242), .B(N220), .S0(N378));
MXI2XL inst_cellmath__53_M_I120 (.Y(inst_cellmath__53_M_out0[10]), .A(N243), .B(N221), .S0(N378));
MXI2XL inst_cellmath__53_M_I121 (.Y(inst_cellmath__53_M_out0[11]), .A(N244), .B(N222), .S0(N378));
MXI2XL inst_cellmath__53_M_I122 (.Y(inst_cellmath__53_M_out0[12]), .A(N245), .B(N223), .S0(N378));
MXI2XL inst_cellmath__53_M_I123 (.Y(inst_cellmath__53_M_out0[13]), .A(N246), .B(N224), .S0(N378));
MXI2XL inst_cellmath__53_M_I124 (.Y(inst_cellmath__53_M_out0[14]), .A(N247), .B(N225), .S0(N378));
MXI2XL inst_cellmath__53_M_I125 (.Y(inst_cellmath__53_M_out0[15]), .A(N248), .B(N226), .S0(N378));
MXI2XL inst_cellmath__53_M_I126 (.Y(inst_cellmath__53_M_out0[16]), .A(N249), .B(N227), .S0(N378));
MXI2XL inst_cellmath__53_M_I127 (.Y(inst_cellmath__53_M_out0[17]), .A(N250), .B(N228), .S0(N378));
MXI2XL inst_cellmath__53_M_I128 (.Y(inst_cellmath__53_M_out0[18]), .A(N251), .B(N229), .S0(N378));
MXI2XL inst_cellmath__53_M_I129 (.Y(inst_cellmath__53_M_out0[19]), .A(N252), .B(N230), .S0(N378));
MXI2XL inst_cellmath__53_M_I130 (.Y(inst_cellmath__53_M_out0[20]), .A(N253), .B(N231), .S0(N378));
MXI2XL inst_cellmath__53_M_I131 (.Y(inst_cellmath__53_M_out0[21]), .A(N254), .B(N232), .S0(N378));
endmodule

/* CADENCE  ubb4SAHWrRw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




