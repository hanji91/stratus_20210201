/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:18 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895;
wire N5143,N5150,N5157,N5164,N5171,N5178,N5185 
	,N5192,N5199,N5206,N5213,N5220,N5227,N5234,N5241 
	,N5248,N5255,N5262,N5269,N5276,N5283,N5295,N5354 
	,N5356,N5592,N5605,N5607,N5631,N5633,N5712,N5717 
	,N5967,N5998,N6004,N6029,N6042,N6048,N6069,N6071 
	,N6079,N6091,N6093,N6099,N6101,N6111,N6119,N6137 
	,N6171,N6182,N6563,N6570,N6572,N6873,N6875,N6880 
	,N6882,N6887,N6889,N6894,N6896,N6899,N6901,N6903 
	,N6908,N6925,N7051,N7053,N7058,N7060,N7063,N7209 
	,N7216,N7318,N7325,N7348,N7368,N7375,N7382,N7389 
	,N7396,N7440,N7536,N7540,N7577,N7604,N7608,N7714 
	,N7720,N7722,N7724,N7727,N7729,N7731,N7998,N8000 
	,N8191,N8192,N8193,N8194;
reg x_reg_15__retimed_I4479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4479_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996;
	end
assign N8000 = x_reg_15__retimed_I4479_QOUT;
reg x_reg_15__retimed_I4478_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4478_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000;
	end
assign N7998 = x_reg_15__retimed_I4478_QOUT;
reg x_reg_15__retimed_I4366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4366_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046;
	end
assign N7731 = x_reg_15__retimed_I4366_QOUT;
reg x_reg_15__retimed_I4365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4365_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061;
	end
assign N7729 = x_reg_15__retimed_I4365_QOUT;
reg x_reg_15__retimed_I4364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4364_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086;
	end
assign N7727 = x_reg_15__retimed_I4364_QOUT;
reg x_reg_15__retimed_I4363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4363_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997;
	end
assign N7724 = x_reg_15__retimed_I4363_QOUT;
reg x_reg_15__retimed_I4362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4362_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070;
	end
assign N7722 = x_reg_15__retimed_I4362_QOUT;
reg x_reg_15__retimed_I4361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4361_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011;
	end
assign N7720 = x_reg_15__retimed_I4361_QOUT;
reg x_reg_15__retimed_I4360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4360_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032;
	end
assign N7714 = x_reg_15__retimed_I4360_QOUT;
reg x_reg_15__retimed_I4344_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4344_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049;
	end
assign N7608 = x_reg_15__retimed_I4344_QOUT;
reg x_reg_15__retimed_I4342_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4342_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078;
	end
assign N7604 = x_reg_15__retimed_I4342_QOUT;
reg x_reg_15__retimed_I4334_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4334_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065;
	end
assign N7577 = x_reg_15__retimed_I4334_QOUT;
reg x_reg_15__retimed_I4331_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4331_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082;
	end
assign N7540 = x_reg_15__retimed_I4331_QOUT;
reg x_reg_15__retimed_I4329_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4329_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014;
	end
assign N7536 = x_reg_15__retimed_I4329_QOUT;
reg x_reg_15__retimed_I4313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4313_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655;
	end
assign N7440 = x_reg_15__retimed_I4313_QOUT;
reg x_reg_15__retimed_I4297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4297_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N7396 = x_reg_15__retimed_I4297_QOUT;
reg x_reg_15__retimed_I4294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4294_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N7389 = x_reg_15__retimed_I4294_QOUT;
reg x_reg_15__retimed_I4291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4291_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N7382 = x_reg_15__retimed_I4291_QOUT;
reg x_reg_15__retimed_I4288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4288_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N7375 = x_reg_15__retimed_I4288_QOUT;
reg x_reg_15__retimed_I4285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4285_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N7368 = x_reg_15__retimed_I4285_QOUT;
reg x_reg_15__retimed_I4277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4277_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N7348 = x_reg_15__retimed_I4277_QOUT;
reg x_reg_15__retimed_I4273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4273_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N7325 = x_reg_15__retimed_I4273_QOUT;
reg x_reg_15__retimed_I4270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4270_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N7318 = x_reg_15__retimed_I4270_QOUT;
reg x_reg_15__retimed_I4238_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4238_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N7216 = x_reg_15__retimed_I4238_QOUT;
reg x_reg_15__retimed_I4235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4235_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N7209 = x_reg_15__retimed_I4235_QOUT;
reg x_reg_15__retimed_I4188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4188_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N7063 = x_reg_15__retimed_I4188_QOUT;
reg x_reg_15__retimed_I4187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4187_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
	end
assign N7060 = x_reg_15__retimed_I4187_QOUT;
reg x_reg_15__retimed_I4186_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4186_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N7058 = x_reg_15__retimed_I4186_QOUT;
reg x_reg_15__retimed_I4184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4184_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18];
	end
assign N7053 = x_reg_15__retimed_I4184_QOUT;
reg x_reg_15__retimed_I4183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4183_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N7051 = x_reg_15__retimed_I4183_QOUT;
reg x_reg_15__retimed_I4139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4139_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N6925 = x_reg_15__retimed_I4139_QOUT;
reg x_reg_15__retimed_I4132_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4132_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N6908 = x_reg_15__retimed_I4132_QOUT;
reg x_reg_15__retimed_I4130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4130_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N6903 = x_reg_15__retimed_I4130_QOUT;
reg x_reg_15__retimed_I4129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4129_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N6901 = x_reg_15__retimed_I4129_QOUT;
reg x_reg_15__retimed_I4128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4128_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N6899 = x_reg_15__retimed_I4128_QOUT;
reg x_reg_15__retimed_I4127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4127_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
	end
assign N6896 = x_reg_15__retimed_I4127_QOUT;
reg x_reg_15__retimed_I4126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4126_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N6894 = x_reg_15__retimed_I4126_QOUT;
reg x_reg_15__retimed_I4124_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4124_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22];
	end
assign N6889 = x_reg_15__retimed_I4124_QOUT;
reg x_reg_15__retimed_I4123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4123_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N6887 = x_reg_15__retimed_I4123_QOUT;
reg x_reg_15__retimed_I4121_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4121_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20];
	end
assign N6882 = x_reg_15__retimed_I4121_QOUT;
reg x_reg_15__retimed_I4120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4120_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N6880 = x_reg_15__retimed_I4120_QOUT;
reg x_reg_15__retimed_I4118_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4118_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19];
	end
assign N6875 = x_reg_15__retimed_I4118_QOUT;
reg x_reg_15__retimed_I4117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4117_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N6873 = x_reg_15__retimed_I4117_QOUT;
reg x_reg_15__retimed_I4000_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I4000_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23];
	end
assign N6572 = x_reg_15__retimed_I4000_QOUT;
reg x_reg_15__retimed_I3999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3999_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15];
	end
assign N6570 = x_reg_15__retimed_I3999_QOUT;
reg x_reg_15__retimed_I3996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3996_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16];
	end
assign N6563 = x_reg_15__retimed_I3996_QOUT;
reg x_reg_15__retimed_I3848_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3848_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N6182 = x_reg_15__retimed_I3848_QOUT;
reg x_reg_15__retimed_I3844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3844_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N6171 = x_reg_15__retimed_I3844_QOUT;
reg x_reg_15__retimed_I3832_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3832_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918;
	end
assign N6137 = x_reg_15__retimed_I3832_QOUT;
reg x_reg_15__retimed_I3825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3825_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944;
	end
assign N6119 = x_reg_15__retimed_I3825_QOUT;
reg x_reg_15__retimed_I3822_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3822_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911;
	end
assign N6111 = x_reg_15__retimed_I3822_QOUT;
reg x_reg_15__retimed_I3818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3818_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923;
	end
assign N6101 = x_reg_15__retimed_I3818_QOUT;
reg x_reg_15__retimed_I3817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3817_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936;
	end
assign N6099 = x_reg_15__retimed_I3817_QOUT;
reg x_reg_15__retimed_I3815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3815_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928;
	end
assign N6093 = x_reg_15__retimed_I3815_QOUT;
reg x_reg_15__retimed_I3814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3814_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N6091 = x_reg_15__retimed_I3814_QOUT;
reg x_reg_15__retimed_I3809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3809_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N6079 = x_reg_15__retimed_I3809_QOUT;
reg x_reg_15__retimed_I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3806_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24];
	end
assign N6071 = x_reg_15__retimed_I3806_QOUT;
reg x_reg_15__retimed_I3805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3805_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
	end
assign N6069 = x_reg_15__retimed_I3805_QOUT;
reg x_reg_15__retimed_I3798_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3798_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901;
	end
assign N6048 = x_reg_15__retimed_I3798_QOUT;
reg x_reg_15__retimed_I3796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3796_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921;
	end
assign N6042 = x_reg_15__retimed_I3796_QOUT;
reg x_reg_15__retimed_I3791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3791_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883;
	end
assign N6029 = x_reg_15__retimed_I3791_QOUT;
reg x_reg_15__retimed_I3783_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3783_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908;
	end
assign N6004 = x_reg_15__retimed_I3783_QOUT;
reg x_reg_15__retimed_I3781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3781_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929;
	end
assign N5998 = x_reg_15__retimed_I3781_QOUT;
reg x_reg_15__retimed_I3768_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3768_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018;
	end
assign N5967 = x_reg_15__retimed_I3768_QOUT;
reg x_reg_23__retimed_I3675_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3675_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N5717 = x_reg_23__retimed_I3675_QOUT;
reg x_reg_22__retimed_I3673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3673_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111;
	end
assign N5712 = x_reg_22__retimed_I3673_QOUT;
reg x_reg_31__retimed_I3668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3668_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N5633 = x_reg_31__retimed_I3668_QOUT;
reg x_reg_31__retimed_I3667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3667_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5631 = x_reg_31__retimed_I3667_QOUT;
reg x_reg_23__retimed_I3659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3659_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5607 = x_reg_23__retimed_I3659_QOUT;
reg x_reg_23__retimed_I3658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3658_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5605 = x_reg_23__retimed_I3658_QOUT;
reg x_reg_15__retimed_I3656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3656_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5592 = x_reg_15__retimed_I3656_QOUT;
assign N8191 = !N5592;
assign N8192 = !N8191;
reg x_reg_31__retimed_I3561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3561_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282;
	end
assign N5356 = x_reg_31__retimed_I3561_QOUT;
reg x_reg_31__retimed_I3560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3560_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291;
	end
assign N5354 = x_reg_31__retimed_I3560_QOUT;
reg x_reg_15__retimed_I3535_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3535_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5295 = x_reg_15__retimed_I3535_QOUT;
reg x_reg_0__retimed_I3530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3530_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5283 = x_reg_0__retimed_I3530_QOUT;
reg x_reg_1__retimed_I3527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3527_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5276 = x_reg_1__retimed_I3527_QOUT;
reg x_reg_2__retimed_I3524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3524_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5269 = x_reg_2__retimed_I3524_QOUT;
reg x_reg_3__retimed_I3521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3521_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5262 = x_reg_3__retimed_I3521_QOUT;
reg x_reg_4__retimed_I3518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3518_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5255 = x_reg_4__retimed_I3518_QOUT;
reg x_reg_5__retimed_I3515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3515_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5248 = x_reg_5__retimed_I3515_QOUT;
reg x_reg_6__retimed_I3512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3512_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5241 = x_reg_6__retimed_I3512_QOUT;
reg x_reg_7__retimed_I3509_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3509_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5234 = x_reg_7__retimed_I3509_QOUT;
reg x_reg_8__retimed_I3506_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3506_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5227 = x_reg_8__retimed_I3506_QOUT;
reg x_reg_9__retimed_I3503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3503_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5220 = x_reg_9__retimed_I3503_QOUT;
reg x_reg_10__retimed_I3500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3500_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5213 = x_reg_10__retimed_I3500_QOUT;
reg x_reg_11__retimed_I3497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3497_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5206 = x_reg_11__retimed_I3497_QOUT;
reg x_reg_12__retimed_I3494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3494_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5199 = x_reg_12__retimed_I3494_QOUT;
reg x_reg_13__retimed_I3491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3491_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5192 = x_reg_13__retimed_I3491_QOUT;
reg x_reg_14__retimed_I3488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3488_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5185 = x_reg_14__retimed_I3488_QOUT;
reg x_reg_16__retimed_I3485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3485_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5178 = x_reg_16__retimed_I3485_QOUT;
reg x_reg_17__retimed_I3482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3482_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5171 = x_reg_17__retimed_I3482_QOUT;
reg x_reg_18__retimed_I3479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3479_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5164 = x_reg_18__retimed_I3479_QOUT;
reg x_reg_19__retimed_I3476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3476_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5157 = x_reg_19__retimed_I3476_QOUT;
reg x_reg_20__retimed_I3473_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3473_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5150 = x_reg_20__retimed_I3473_QOUT;
reg x_reg_21__retimed_I3470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3470_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5143 = x_reg_21__retimed_I3470_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4132 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8834);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172 = !(((a_man[0] | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4168);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4174) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4163) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4183);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4172) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4166) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4177) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4187);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221 = !(((b_exp[5] & b_exp[4]) & b_exp[7]) & b_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218 = !(((b_exp[0] & b_exp[1]) & b_exp[2]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4221 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4218);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4245);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4232 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4251) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4240) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4260);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4249) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4243) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4254) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4264);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408 = a_exp[7] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 = a_exp[6] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 = a_exp[5] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 = a_exp[4] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 = a_exp[3] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 = a_exp[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733 = !a_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8733) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557) & a_exp[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8730;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404 = !(a_exp[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372 = a_exp[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380 = !(a_exp[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8840) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377 = a_exp[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417 = a_exp[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382 = a_exp[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357 = a_exp[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393 = !(a_exp[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 | a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4380;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8847) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4377) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4417) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4382) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4357) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4393;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8854) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607 = !a_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489 = !(b_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542 = !(b_man[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4542);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4568);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473 = !a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 = !(b_man[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496 = !(b_man[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4496);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548 = !(b_man[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600 = !(b_man[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4550 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552 = !a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559 = !(b_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613 = !(b_man[10] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4613);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514 = !(b_man[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516 = !a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502 = !(b_man[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555 = !(b_man[14] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4555);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605 = !(b_man[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509 = !(b_man[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4509);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4530);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566 = !(b_man[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4566);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588 = !a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467 = !(b_man[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518 = !(b_man[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4518);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610 = !a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569 = !(b_man[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471 = !(b_man[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4471);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4491);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523 = !(b_man[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4497);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590 = !(((a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4504) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4477) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4512);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4523)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4590 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4558) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4543);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4506) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4569)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4524);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4588);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4551) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4467)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4500);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4611 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4576) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4545);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4599) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4567)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4533);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4570);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4514)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4546);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4484);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4552);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4493) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4559)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4591);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4479 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4565);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4531);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4540) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4605)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4487);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4598);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4516);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4587) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4502)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4534);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4499 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4466) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4469) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4553);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4495 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4614) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4580);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4482) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4548)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4581);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4561);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4473);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4528) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4476);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4517 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4483) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4602);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4541);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4607);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4574) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4489)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4522);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4536 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4538) | (b_man[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4520));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4486) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4571));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4562) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4510)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4475);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[8] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4310 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4314);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340 = ((b_exp[7] | b_exp[5]) | b_exp[6]) | b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336 = ((b_exp[0] | b_exp[1]) | b_exp[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4340 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4336);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4414 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4375) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4408;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4407 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4384) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4396;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4368 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4404) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4364;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8738 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4402 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4387) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4386;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4390 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4405) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4379 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4370) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4376;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4373 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4401) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4418;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4793) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4792 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8749;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = a_exp[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 = a_exp[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4751) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4989 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5023 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5107 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5110 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5059 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5062));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5010 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5013 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8882;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4921 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5100 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4958 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5070 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8875;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4995 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4998 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5097 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5120 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8868;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4939 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & a_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8861;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5084 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5061));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4930);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5012 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5021);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5096);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4969));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4929);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4955);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5089 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5047);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5103);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5068);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4946);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4976);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5048);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5104));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4915);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4991 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5075);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4984);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4954);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5428 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5400);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5008 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4906);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5028);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5055 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4982);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5095);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5002);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5000 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5411);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5414);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5027) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5085 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4923);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5015);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5112);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5398 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5408);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5419 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5082 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5416 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5427 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5397);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5418 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5436;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N625 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8708;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5767);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N656 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N657 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5742);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5792)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5749);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N659 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N660 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5695);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5766)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5723);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5771) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5728);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5672);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5644);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5741)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5702);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5791);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5717)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5679);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5745) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5698)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5655);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5684 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5687) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5831;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5664;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5816;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5827)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5674);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5785;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5811) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5659);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5819)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5837;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5701 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5714;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5730;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5756)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5800);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5646) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5665;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5840 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5772;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5660)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5813);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5753);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5781 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5689;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5838) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5798;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5051);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4960);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4990);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5111);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5014);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & a_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5342) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4953) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4922);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5465;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5721);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5682 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5809) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5765);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5694)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5651);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5737 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5836) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5790);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5715);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5693);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5823));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5671) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5775 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5822) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5778)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5801);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5803 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5731;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5650) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5648;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5691;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5830 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5758;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5675;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5750) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5805)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5656);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5657 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5783;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5677) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5700;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010 = !(N7720 & N7729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5686;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5839;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5773) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5820);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5806;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5744)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5835) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5735;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5661;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5710)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5752);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5796) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5786;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5668 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5703;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5832);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5770 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5760;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5643) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5680;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5763;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5779);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5808 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5711;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5793) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5824;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6065 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6073);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6083 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6063));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6019;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6009 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5998) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6028);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6047 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6026));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6076;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6078 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6054) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031 = !((N7608 & N7729) | N7604);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] = ((!N7577) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6031);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919 = (!N6171) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6033);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6006);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5725) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5814;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6038) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6057);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6067) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6087);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6079) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6015);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6032 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6004);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6001) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6021);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6029) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6050);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6046 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6043) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6071);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6058) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6080);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5993) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6016);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6086 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6007) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6035);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074 = !((N7731 & N7729) | N7727);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0] = ((!N7714) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6074);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6014 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6041 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6060));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6069));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6024;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6082 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6042) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6005)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6062);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010) & (!N7536)) | (!N7540));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0];
assign N8193 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416;
assign N8194 = !N8193;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039 = !(N7998 & N8000);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6000 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5996));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6061;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439 = (N7720 & N7722) | N7724;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 & N7389;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6882) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6880);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6328 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 & N7396;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6875) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6873);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6457 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6416;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8804;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7216) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7368);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6071) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6563);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6307 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7209;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6572) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6570);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6436 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6423 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6367 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809 & N7375;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N7053) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N7051);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6420 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383 = N7382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8809;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N7060) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N7058);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6386 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7318;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6889) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6887);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6400 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7325;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6896) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N6894);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6365 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6459 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6326 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6408 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6389 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6352 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6330 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439 & N7368;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6563) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N7216);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6347) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6349 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6337 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6318 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6444 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6422 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6453 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N6887) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7318);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6441 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N6894) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7325);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6405 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6317 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N6880) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7389);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N6873) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7396);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6334 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806 & N6570) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8806) & N7209);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6315 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6300 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6414 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6344 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6443 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7051) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7375);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6297 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6435 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6395 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6324 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6373 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6402 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6407 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6387 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6438 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808 & N7058) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8808) & N7382);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6427 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6364 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6335 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6321 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6429 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6456 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6385 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6298 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6411 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6314 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6394 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6331 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6424 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6368 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6341 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6404 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6357 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6361 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8812;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6448 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6333 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6426 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6323 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6454);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6355 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6390 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6319 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6353 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6445 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6383);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6447 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6312);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6452 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6306 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6434 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6377 & N8194) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6303 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8814));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6343) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6397 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6301 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6375));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6409 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6338 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6362 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N6908) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 & a_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32) & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6398);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6419 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8772;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6655 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6308) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1])) | (!N7440);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N7348) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633 = N7063 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636 = !(((N6903 | N6901) | N6899) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639 = !(N6925 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N636) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__53)) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6430 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6450 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6358 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8824) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6380 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6749 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6417 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6346 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8820) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6310 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6775);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951 = N6182 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941 = !(N6182 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6941);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909 = !(N6171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6909);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[2]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6918} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946 = N6137 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N2691) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[3]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6944} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6931};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913 = (!N6119) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6946) | (!(N6137 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6360)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917)) | ((!N6119) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6439));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[4]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6911} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6902};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938 = N6111 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6938) | (!(N6111 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6311)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6908 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6936) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6923;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932) ^ N6004;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905 = ((!N6004) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6932)) | ((!N6099) & (!N6101));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6929 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6928;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905) ^ N5998;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6905 & N5998) | (!(N6091 | N6093)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6901 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6921;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930) ^ N6048;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950 = ((!N6048) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6930)) | ((!N6079) & (!N6042));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = (!N6042) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6951;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6948) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6919;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6917) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6913;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6999);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7018 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6010 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6039);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6883 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6889));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] & N6071) | N6069);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62 = !(N6029 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = N6042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020 = !(((N5967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7000) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8722)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7020));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074 | (!N8192));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7092);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7111 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70 = N5712 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 = !(N8192 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8825;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6720) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7182 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6777 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7138) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5143);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6703;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6714) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7195) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5150);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6721 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7153) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5157);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6768;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6767 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6705) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8826 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7207) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5164);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8830;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13892;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6766 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7166) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5171);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6732;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6696) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7122) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5178);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6702 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5295);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6751 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6727 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6770) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7133) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5185);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6758 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7190) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5192);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6695;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6729) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7146) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5199);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6762 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7202) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5206);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6709 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6763) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7161) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5213);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6718 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7117) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5220);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6759;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6754) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7173) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5227);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6744 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7129) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5234);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6719 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6748) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7186) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5241);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6713 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7142) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5248);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6710) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7198) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5255);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6731 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7156) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5262);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6701 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7210) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5269);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6776) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7169) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5276);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[0]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7150 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13893 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7125) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7141 & N5283);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068 = ((N5605 | N5607) | N5592) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7074;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7068) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651 = N5717 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0] = ((N5605 | N5607) | N8192) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N7056) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8785);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13895 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6212 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6233);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6282 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] & N5633) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]) & N5631);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6291 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706);
assign x[31] = (N5354 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6285) | ((!N5354) & N5356);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__28[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLbzSg7aoxA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



