/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:24 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_3_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417;
wire N8340,N8378,N8385,N8392,N8398,N8401,N8410 
	,N8419,N8428,N8437,N8446,N8455,N8464,N8473,N8482 
	,N8491,N8500,N8509,N8518,N8527,N8536,N8545,N8554 
	,N8563,N8572,N8581,N8790,N8795,N8800,N8805,N8810 
	,N8815,N8820,N8825,N8830,N8835,N8840,N8845,N8850 
	,N8855,N8860,N8865,N8870,N8875,N8880,N8885,N8890 
	,N8895,N8939,N8965,N8991,N9320,N9322,N9377,N9379 
	,N9386,N9388,N9395,N9397,N9404,N9406,N9413,N9415 
	,N9422,N9424,N9431,N9433,N9440,N9442,N9449,N9451 
	,N9457,N9459,N9500,N9502,N9504,N9518,N9520,N9545 
	,N9808,N9814,N9820,N9826,N9832,N9838,N9844,N9850 
	,N9872,N9874,N9892,N9894,N9902,N9912,N9914,N9922 
	,N9924,N9932,N9934,N10016,N10018,N10023,N10025,N10030 
	,N10032,N10037,N10039,N10046,N10051,N10058,N10060,N10065 
	,N10074,N10079,N10081,N10100,N10102,N10107,N10121,N10123 
	,N10128,N10153,N10159,N10163,N10165,N10169,N10171,N10274 
	,N10277,N10285,N10293,N10301,N10309,N10317,N10325,N10333 
	,N10341,N10349,N10357,N10995,N10996;
reg x_reg_21__retimed_I5666_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5666_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501;
	end
assign N10357 = x_reg_21__retimed_I5666_QOUT;
reg x_reg_21__retimed_I5663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5663_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320;
	end
assign N10349 = x_reg_21__retimed_I5663_QOUT;
reg x_reg_21__retimed_I5660_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5660_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591;
	end
assign N10341 = x_reg_21__retimed_I5660_QOUT;
reg x_reg_21__retimed_I5657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5657_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407;
	end
assign N10333 = x_reg_21__retimed_I5657_QOUT;
reg x_reg_21__retimed_I5654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5654_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672;
	end
assign N10325 = x_reg_21__retimed_I5654_QOUT;
reg x_reg_21__retimed_I5651_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5651_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475;
	end
assign N10317 = x_reg_21__retimed_I5651_QOUT;
reg x_reg_21__retimed_I5648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5648_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755;
	end
assign N10309 = x_reg_21__retimed_I5648_QOUT;
reg x_reg_21__retimed_I5645_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5645_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561;
	end
assign N10301 = x_reg_21__retimed_I5645_QOUT;
reg x_reg_21__retimed_I5642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5642_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840;
	end
assign N10293 = x_reg_21__retimed_I5642_QOUT;
reg x_reg_21__retimed_I5639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5639_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645;
	end
assign N10285 = x_reg_21__retimed_I5639_QOUT;
reg x_reg_21__retimed_I5636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5636_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917;
	end
assign N10277 = x_reg_21__retimed_I5636_QOUT;
reg x_reg_21__retimed_I5635_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5635_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178;
	end
assign N10274 = x_reg_21__retimed_I5635_QOUT;
reg x_reg_21__retimed_I5613_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5613_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821;
	end
assign N10171 = x_reg_21__retimed_I5613_QOUT;
reg x_reg_21__retimed_I5612_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5612_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310;
	end
assign N10169 = x_reg_21__retimed_I5612_QOUT;
reg x_reg_21__retimed_I5611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5611_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483;
	end
assign N10165 = x_reg_21__retimed_I5611_QOUT;
reg x_reg_21__retimed_I5610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5610_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081;
	end
assign N10163 = x_reg_21__retimed_I5610_QOUT;
reg x_reg_21__retimed_I5609_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5609_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617;
	end
assign N10159 = x_reg_21__retimed_I5609_QOUT;
reg x_reg_21__retimed_I5607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5607_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293;
	end
assign N10153 = x_reg_21__retimed_I5607_QOUT;
reg x_reg_21__retimed_I5597_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5597_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0];
	end
assign N10128 = x_reg_21__retimed_I5597_QOUT;
reg x_reg_21__retimed_I5595_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5595_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18];
	end
assign N10123 = x_reg_21__retimed_I5595_QOUT;
reg x_reg_21__retimed_I5594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5594_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17];
	end
assign N10121 = x_reg_21__retimed_I5594_QOUT;
reg x_reg_21__retimed_I5588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5588_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19];
	end
assign N10107 = x_reg_21__retimed_I5588_QOUT;
reg x_reg_21__retimed_I5586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5586_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21];
	end
assign N10102 = x_reg_21__retimed_I5586_QOUT;
reg x_reg_21__retimed_I5585_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5585_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20];
	end
assign N10100 = x_reg_21__retimed_I5585_QOUT;
reg x_reg_21__retimed_I5577_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5577_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12];
	end
assign N10081 = x_reg_21__retimed_I5577_QOUT;
reg x_reg_21__retimed_I5576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5576_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11];
	end
assign N10079 = x_reg_21__retimed_I5576_QOUT;
reg x_reg_21__retimed_I5574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5574_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7];
	end
assign N10074 = x_reg_21__retimed_I5574_QOUT;
reg x_reg_21__retimed_I5570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5570_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3];
	end
assign N10065 = x_reg_21__retimed_I5570_QOUT;
reg x_reg_21__retimed_I5568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5568_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14];
	end
assign N10060 = x_reg_21__retimed_I5568_QOUT;
reg x_reg_21__retimed_I5567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5567_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13];
	end
assign N10058 = x_reg_21__retimed_I5567_QOUT;
reg x_reg_21__retimed_I5564_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5564_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8];
	end
assign N10051 = x_reg_21__retimed_I5564_QOUT;
reg x_reg_21__retimed_I5562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5562_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6];
	end
assign N10046 = x_reg_21__retimed_I5562_QOUT;
reg x_reg_21__retimed_I5559_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5559_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10];
	end
assign N10039 = x_reg_21__retimed_I5559_QOUT;
reg x_reg_21__retimed_I5558_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5558_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9];
	end
assign N10037 = x_reg_21__retimed_I5558_QOUT;
reg x_reg_21__retimed_I5556_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5556_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5];
	end
assign N10032 = x_reg_21__retimed_I5556_QOUT;
reg x_reg_21__retimed_I5555_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5555_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4];
	end
assign N10030 = x_reg_21__retimed_I5555_QOUT;
reg x_reg_21__retimed_I5553_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5553_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2];
	end
assign N10025 = x_reg_21__retimed_I5553_QOUT;
reg x_reg_21__retimed_I5552_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5552_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1];
	end
assign N10023 = x_reg_21__retimed_I5552_QOUT;
reg x_reg_21__retimed_I5550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5550_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16];
	end
assign N10018 = x_reg_21__retimed_I5550_QOUT;
reg x_reg_21__retimed_I5549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5549_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15];
	end
assign N10016 = x_reg_21__retimed_I5549_QOUT;
reg x_reg_21__retimed_I5521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5521_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33];
	end
assign N9934 = x_reg_21__retimed_I5521_QOUT;
reg x_reg_21__retimed_I5520_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5520_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32];
	end
assign N9932 = x_reg_21__retimed_I5520_QOUT;
reg x_reg_21__retimed_I5518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5518_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31];
	end
assign N9924 = x_reg_21__retimed_I5518_QOUT;
reg x_reg_21__retimed_I5517_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5517_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30];
	end
assign N9922 = x_reg_21__retimed_I5517_QOUT;
reg x_reg_21__retimed_I5515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5515_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25];
	end
assign N9914 = x_reg_21__retimed_I5515_QOUT;
reg x_reg_21__retimed_I5514_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5514_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24];
	end
assign N9912 = x_reg_21__retimed_I5514_QOUT;
reg x_reg_21__retimed_I5511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5511_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34];
	end
assign N9902 = x_reg_21__retimed_I5511_QOUT;
reg x_reg_21__retimed_I5509_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5509_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29];
	end
assign N9894 = x_reg_21__retimed_I5509_QOUT;
reg x_reg_21__retimed_I5508_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5508_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28];
	end
assign N9892 = x_reg_21__retimed_I5508_QOUT;
reg x_reg_21__retimed_I5503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5503_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27];
	end
assign N9874 = x_reg_21__retimed_I5503_QOUT;
reg x_reg_21__retimed_I5502_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5502_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26];
	end
assign N9872 = x_reg_21__retimed_I5502_QOUT;
reg x_reg_21__retimed_I5494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5494_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415;
	end
assign N9850 = x_reg_21__retimed_I5494_QOUT;
reg x_reg_21__retimed_I5492_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5492_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100;
	end
assign N9844 = x_reg_21__retimed_I5492_QOUT;
reg x_reg_21__retimed_I5490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5490_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219;
	end
assign N9838 = x_reg_21__retimed_I5490_QOUT;
reg x_reg_21__retimed_I5488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5488_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900;
	end
assign N9832 = x_reg_21__retimed_I5488_QOUT;
reg x_reg_21__retimed_I5486_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5486_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571;
	end
assign N9826 = x_reg_21__retimed_I5486_QOUT;
reg x_reg_21__retimed_I5484_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5484_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704;
	end
assign N9820 = x_reg_21__retimed_I5484_QOUT;
reg x_reg_21__retimed_I5482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5482_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379;
	end
assign N9814 = x_reg_21__retimed_I5482_QOUT;
reg x_reg_21__retimed_I5480_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5480_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503;
	end
assign N9808 = x_reg_21__retimed_I5480_QOUT;
reg x_reg_21__retimed_I5394_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5394_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4;
	end
assign N9545 = x_reg_21__retimed_I5394_QOUT;
reg x_reg_21__retimed_I5387_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5387_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23];
	end
assign N9520 = x_reg_21__retimed_I5387_QOUT;
reg x_reg_21__retimed_I5386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5386_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22];
	end
assign N9518 = x_reg_21__retimed_I5386_QOUT;
reg x_reg_21__retimed_I5380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5380_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446;
	end
assign N9504 = x_reg_21__retimed_I5380_QOUT;
reg x_reg_21__retimed_I5379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5379_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445;
	end
assign N9502 = x_reg_21__retimed_I5379_QOUT;
reg x_reg_21__retimed_I5378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5378_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8;
	end
assign N9500 = x_reg_21__retimed_I5378_QOUT;
reg x_reg_21__retimed_I5366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5366_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8];
	end
assign N9459 = x_reg_21__retimed_I5366_QOUT;
reg x_reg_21__retimed_I5365_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5365_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8];
	end
assign N9457 = x_reg_21__retimed_I5365_QOUT;
reg x_reg_21__retimed_I5363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5363_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1];
	end
assign N9451 = x_reg_21__retimed_I5363_QOUT;
reg x_reg_21__retimed_I5362_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5362_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1];
	end
assign N9449 = x_reg_21__retimed_I5362_QOUT;
reg x_reg_21__retimed_I5360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5360_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3];
	end
assign N9442 = x_reg_21__retimed_I5360_QOUT;
reg x_reg_21__retimed_I5359_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5359_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3];
	end
assign N9440 = x_reg_21__retimed_I5359_QOUT;
reg x_reg_21__retimed_I5357_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5357_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6];
	end
assign N9433 = x_reg_21__retimed_I5357_QOUT;
reg x_reg_21__retimed_I5356_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5356_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6];
	end
assign N9431 = x_reg_21__retimed_I5356_QOUT;
reg x_reg_21__retimed_I5354_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5354_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
	end
assign N9424 = x_reg_21__retimed_I5354_QOUT;
reg x_reg_21__retimed_I5353_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5353_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7];
	end
assign N9422 = x_reg_21__retimed_I5353_QOUT;
reg x_reg_21__retimed_I5351_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5351_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9];
	end
assign N9415 = x_reg_21__retimed_I5351_QOUT;
reg x_reg_21__retimed_I5350_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5350_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9];
	end
assign N9413 = x_reg_21__retimed_I5350_QOUT;
reg x_reg_21__retimed_I5348_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5348_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5];
	end
assign N9406 = x_reg_21__retimed_I5348_QOUT;
reg x_reg_21__retimed_I5347_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5347_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5];
	end
assign N9404 = x_reg_21__retimed_I5347_QOUT;
reg x_reg_21__retimed_I5345_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5345_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4];
	end
assign N9397 = x_reg_21__retimed_I5345_QOUT;
reg x_reg_21__retimed_I5344_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5344_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4];
	end
assign N9395 = x_reg_21__retimed_I5344_QOUT;
reg x_reg_21__retimed_I5342_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5342_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2];
	end
assign N9388 = x_reg_21__retimed_I5342_QOUT;
reg x_reg_21__retimed_I5341_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5341_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2];
	end
assign N9386 = x_reg_21__retimed_I5341_QOUT;
reg x_reg_21__retimed_I5339_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5339_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0];
	end
assign N9379 = x_reg_21__retimed_I5339_QOUT;
reg x_reg_21__retimed_I5338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5338_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0];
	end
assign N9377 = x_reg_21__retimed_I5338_QOUT;
reg x_reg_21__retimed_I5316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5316_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27;
	end
assign N9322 = x_reg_21__retimed_I5316_QOUT;
reg x_reg_21__retimed_I5315_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5315_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28;
	end
assign N9320 = x_reg_21__retimed_I5315_QOUT;
reg x_reg_21__retimed_I5200_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5200_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26;
	end
assign N8991 = x_reg_21__retimed_I5200_QOUT;
reg x_reg_21__retimed_I5198_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5198_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014;
	end
assign N8965 = x_reg_21__retimed_I5198_QOUT;
reg x_reg_21__retimed_I5196_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5196_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095;
	end
assign N8939 = x_reg_21__retimed_I5196_QOUT;
reg x_reg_21__retimed_I5190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5190_QOUT <= a_man[21];
	end
assign N8895 = x_reg_21__retimed_I5190_QOUT;
reg x_reg_20__retimed_I5188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I5188_QOUT <= a_man[20];
	end
assign N8890 = x_reg_20__retimed_I5188_QOUT;
reg x_reg_19__retimed_I5186_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I5186_QOUT <= a_man[19];
	end
assign N8885 = x_reg_19__retimed_I5186_QOUT;
reg x_reg_18__retimed_I5184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I5184_QOUT <= a_man[18];
	end
assign N8880 = x_reg_18__retimed_I5184_QOUT;
reg x_reg_17__retimed_I5182_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I5182_QOUT <= a_man[17];
	end
assign N8875 = x_reg_17__retimed_I5182_QOUT;
reg x_reg_16__retimed_I5180_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I5180_QOUT <= a_man[16];
	end
assign N8870 = x_reg_16__retimed_I5180_QOUT;
reg x_reg_15__retimed_I5178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I5178_QOUT <= a_man[15];
	end
assign N8865 = x_reg_15__retimed_I5178_QOUT;
reg x_reg_14__retimed_I5176_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I5176_QOUT <= a_man[14];
	end
assign N8860 = x_reg_14__retimed_I5176_QOUT;
reg x_reg_13__retimed_I5174_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I5174_QOUT <= a_man[13];
	end
assign N8855 = x_reg_13__retimed_I5174_QOUT;
reg x_reg_12__retimed_I5172_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I5172_QOUT <= a_man[12];
	end
assign N8850 = x_reg_12__retimed_I5172_QOUT;
reg x_reg_11__retimed_I5170_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I5170_QOUT <= a_man[11];
	end
assign N8845 = x_reg_11__retimed_I5170_QOUT;
reg x_reg_10__retimed_I5168_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I5168_QOUT <= a_man[10];
	end
assign N8840 = x_reg_10__retimed_I5168_QOUT;
reg x_reg_9__retimed_I5166_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I5166_QOUT <= a_man[9];
	end
assign N8835 = x_reg_9__retimed_I5166_QOUT;
reg x_reg_8__retimed_I5164_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I5164_QOUT <= a_man[8];
	end
assign N8830 = x_reg_8__retimed_I5164_QOUT;
reg x_reg_7__retimed_I5162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I5162_QOUT <= a_man[7];
	end
assign N8825 = x_reg_7__retimed_I5162_QOUT;
reg x_reg_6__retimed_I5160_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I5160_QOUT <= a_man[6];
	end
assign N8820 = x_reg_6__retimed_I5160_QOUT;
reg x_reg_5__retimed_I5158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I5158_QOUT <= a_man[5];
	end
assign N8815 = x_reg_5__retimed_I5158_QOUT;
reg x_reg_4__retimed_I5156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I5156_QOUT <= a_man[4];
	end
assign N8810 = x_reg_4__retimed_I5156_QOUT;
reg x_reg_3__retimed_I5154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I5154_QOUT <= a_man[3];
	end
assign N8805 = x_reg_3__retimed_I5154_QOUT;
reg x_reg_2__retimed_I5152_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I5152_QOUT <= a_man[2];
	end
assign N8800 = x_reg_2__retimed_I5152_QOUT;
reg x_reg_1__retimed_I5150_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I5150_QOUT <= a_man[1];
	end
assign N8795 = x_reg_1__retimed_I5150_QOUT;
reg x_reg_0__retimed_I5148_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I5148_QOUT <= a_man[0];
	end
assign N8790 = x_reg_0__retimed_I5148_QOUT;
reg x_reg_21__retimed_I5055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5055_QOUT <= b_man[21];
	end
assign N8581 = x_reg_21__retimed_I5055_QOUT;
reg x_reg_20__retimed_I5051_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I5051_QOUT <= b_man[20];
	end
assign N8572 = x_reg_20__retimed_I5051_QOUT;
reg x_reg_19__retimed_I5047_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I5047_QOUT <= b_man[19];
	end
assign N8563 = x_reg_19__retimed_I5047_QOUT;
reg x_reg_18__retimed_I5043_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I5043_QOUT <= b_man[18];
	end
assign N8554 = x_reg_18__retimed_I5043_QOUT;
reg x_reg_17__retimed_I5039_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I5039_QOUT <= b_man[17];
	end
assign N8545 = x_reg_17__retimed_I5039_QOUT;
reg x_reg_16__retimed_I5035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I5035_QOUT <= b_man[16];
	end
assign N8536 = x_reg_16__retimed_I5035_QOUT;
reg x_reg_15__retimed_I5031_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I5031_QOUT <= b_man[15];
	end
assign N8527 = x_reg_15__retimed_I5031_QOUT;
reg x_reg_14__retimed_I5027_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I5027_QOUT <= b_man[14];
	end
assign N8518 = x_reg_14__retimed_I5027_QOUT;
reg x_reg_13__retimed_I5023_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I5023_QOUT <= b_man[13];
	end
assign N8509 = x_reg_13__retimed_I5023_QOUT;
reg x_reg_12__retimed_I5019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I5019_QOUT <= b_man[12];
	end
assign N8500 = x_reg_12__retimed_I5019_QOUT;
reg x_reg_11__retimed_I5015_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I5015_QOUT <= b_man[11];
	end
assign N8491 = x_reg_11__retimed_I5015_QOUT;
reg x_reg_10__retimed_I5011_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I5011_QOUT <= b_man[10];
	end
assign N8482 = x_reg_10__retimed_I5011_QOUT;
reg x_reg_9__retimed_I5007_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I5007_QOUT <= b_man[9];
	end
assign N8473 = x_reg_9__retimed_I5007_QOUT;
reg x_reg_8__retimed_I5003_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I5003_QOUT <= b_man[8];
	end
assign N8464 = x_reg_8__retimed_I5003_QOUT;
reg x_reg_7__retimed_I4999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I4999_QOUT <= b_man[7];
	end
assign N8455 = x_reg_7__retimed_I4999_QOUT;
reg x_reg_6__retimed_I4995_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I4995_QOUT <= b_man[6];
	end
assign N8446 = x_reg_6__retimed_I4995_QOUT;
reg x_reg_5__retimed_I4991_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I4991_QOUT <= b_man[5];
	end
assign N8437 = x_reg_5__retimed_I4991_QOUT;
reg x_reg_4__retimed_I4987_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I4987_QOUT <= b_man[4];
	end
assign N8428 = x_reg_4__retimed_I4987_QOUT;
reg x_reg_3__retimed_I4983_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I4983_QOUT <= b_man[3];
	end
assign N8419 = x_reg_3__retimed_I4983_QOUT;
reg x_reg_2__retimed_I4979_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I4979_QOUT <= b_man[2];
	end
assign N8410 = x_reg_2__retimed_I4979_QOUT;
reg x_reg_1__retimed_I4975_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I4975_QOUT <= b_man[1];
	end
assign N8401 = x_reg_1__retimed_I4975_QOUT;
reg x_reg_0__retimed_I4974_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I4974_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47;
	end
assign N8398 = x_reg_0__retimed_I4974_QOUT;
assign N10995 = !N8398;
assign N10996 = !N10995;
reg x_reg_0__retimed_I4971_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I4971_QOUT <= b_man[0];
	end
assign N8392 = x_reg_0__retimed_I4971_QOUT;
reg x_reg_22__retimed_I4968_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4968_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925;
	end
assign N8385 = x_reg_22__retimed_I4968_QOUT;
reg x_reg_23__retimed_I4965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I4965_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893;
	end
assign N8378 = x_reg_23__retimed_I4965_QOUT;
reg x_reg_29__retimed_I4949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I4949_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874;
	end
assign N8340 = x_reg_29__retimed_I4949_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011 = !(a_exp[0] & a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396 = !((a_exp[7] & a_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900 = !(b_exp[0] & b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388 = !((b_exp[7] & b_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940 = !(((b_man[0] | b_man[1]) | b_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923 = !(b_man[10] | b_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942 = !(b_man[6] | b_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931 = !(b_man[8] | b_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951 = !(b_man[4] | b_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096 = !(b_exp[0] | b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103 = !(b_exp[5] | b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100 = !(b_exp[7] | b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091 = !(b_exp[3] | b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0] = (!b_exp[0]) ^ a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134 = !a_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320 = (!b_man[22]) ^ b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452 = !a_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799 = !a_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963 = b_man[22] | b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385 = (!b_man[20]) ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118 = b_man[21] ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395 = !b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329 = !a_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660 = !a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450 = (!b_man[18]) ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325 = b_man[19] ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993 = !b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653 = !a_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987 = !a_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090 = b_man[17] ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519 = (!b_man[16]) ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583 = !b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513 = !a_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308 = !a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586 = (!b_man[14]) ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295 = b_man[15] ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352 = !b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853 = !a_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186 = !a_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646 = (!b_man[12]) ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060 = b_man[13] ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947 = !b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171 = !a_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511 = !a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712 = (!b_man[10]) ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267 = b_man[11] ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258 = !b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047 = !a_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391 = !a_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779 = (!b_man[8]) ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033 = b_man[9] ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564 = !b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368 = !a_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713 = !a_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844 = (!b_man[6]) ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242 = b_man[7] ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332 = !b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243 = !a_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578 = !a_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906 = b_man[4] ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004 = (!b_man[5]) ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645 = !b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573 = !a_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911 = !a_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968 = (!b_man[2]) ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211 = b_man[3] ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959 = !b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228 = !a_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445 = !a_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272 = !b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357 = !b_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807 = !(b_man[21] & b_man[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529 = !(b_man[19] & b_man[20]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871 = b_man[21] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595 = !(b_man[17] & b_man[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933 = b_man[19] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658 = !(b_man[15] & b_man[16]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994 = b_man[17] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721 = !(b_man[13] & b_man[14]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058 = b_man[15] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795 = !(b_man[11] & b_man[12]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126 = b_man[13] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855 = !(b_man[9] & b_man[10]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185 = b_man[11] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916 = !(b_man[7] & b_man[8]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251 = b_man[9] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978 = !(b_man[5] & b_man[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317 = b_man[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045 = !(b_man[3] & b_man[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385 = b_man[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111 = !(b_man[1] & b_man[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446 = b_man[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435 = b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558) & (!(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922) & (!(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516 = (!N10357) | (N10163 & N10165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104 = (!N10349) | (N10159 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349 = (!N10341) | (N10153 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723 = (!N10333) | (N9850 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776 = (!N10325) | (N9844 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493 = (!N10317) | (N9838 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356 = (!N10309) | (N9832 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331 = (!N10301) | (N9826 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526 = (!N10293) | (N9820 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315 = (!N10285) | (N9814 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326 = (!N10277) | (N9808 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326 ^ N10274;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315) ^ N9808;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356) ^ N9826;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331) ^ N9820;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493) ^ N9832;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526) ^ N9814;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9922) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9894);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9894) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9892);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9892) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9874);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9874) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9872);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9872) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9914);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9914) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9912);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9912) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9520);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516) ^ N10159;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104) ^ N10153;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36] = (!N10163) ^ N10165;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35] = (!N10169) ^ N10171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9902);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9902) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9934) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9932);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9932) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9924);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9924) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9922);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776) ^ N9838;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723) ^ N9844;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349) ^ N9850;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9520) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N9518);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23 = a_sign ^ b_sign;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10039) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10037);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10060) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10058);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10081) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10079);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10018) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10016);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10025) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10023);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10046) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10032);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10030) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10065);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10051) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10074);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10032) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10030);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10037) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10051);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10074) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10046);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10079) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10039);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10065) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10025);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N9518) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10102);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10100) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10107);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10123) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10121);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0] = b_man[1] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10128;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N10023) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N10128);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10102) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10100);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N10107) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N10123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N10121) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N10018);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N10016) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N10060);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N10058) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N10081);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24])) | (!N9545));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447 = ((N9500 | N9502) | N9504) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450 = ((!N9504) & (!N9502)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9379) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631 = b_exp[0] | a_exp[0];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]} = {1'B0, a_exp[1]} + {1'B0, b_exp[1]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]} = {1'B0, a_exp[2]} + {1'B0, b_exp[2]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9388) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9386);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]} = {1'B0, a_exp[3]} + {1'B0, b_exp[3]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]} = {1'B0, a_exp[4]} + {1'B0, b_exp[4]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9397) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9395);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]} = {1'B0, a_exp[5]} + {1'B0, b_exp[5]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9406) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9404);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5]);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]} = {1'B0, a_exp[6]} + {1'B0, b_exp[6]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627 = !a_exp[7];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]} = {1'B0, b_exp[7]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9424) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9422);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9442) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9440);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] = (!a_exp[7]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9459) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9457);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9451) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9449);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9433) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9431);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9] = !(a_exp[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N9415) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N9413);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830 = !(((N9320 | N9322) | N8991) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 = !(N8939 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8895);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 = !(N8965 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 = !(N8991 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852 = !(rm[0] & rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7 = !(rm[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8581) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[21] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8890);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8572) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[20] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8885);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8563) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[19] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8880);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8554) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[18] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8875);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8545) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[17] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8870);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8536) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[16] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8865);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8527) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[15] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8860);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8518) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[14] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8855);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8509) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[13] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8850);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8500) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[12] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8491) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[11] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8840);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8482) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[10] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8835);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8473) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[9] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8830);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8464) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[8] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8825);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8455) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8820);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8446) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8815);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8437) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[5] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8810);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8428) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8805);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8419) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[3] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8800);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8410) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[2] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8795);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8401) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[1] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N8790);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 & N8392) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N10996));
assign x[0] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47);
assign x[22] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49 & N8385) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887;
assign x[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7]);
assign x[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6]);
assign x[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5]);
assign x[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4]);
assign x[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3]);
assign x[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2]);
assign x[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8340) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470);
assign x[23] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N8378) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 & (!b_sign));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 & a_sign) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23);
reg x_reg_31__I1625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I1625_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31];
	end
assign x[31] = x_reg_31__I1625_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vrj1TwrfrB4= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



