/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:38:04 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_5_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
wire N5507,N5514,N5521,N5528,N5535,N5542,N5549 
	,N5556,N5563,N5570,N5577,N5584,N5591,N5598,N5605 
	,N5612,N5619,N5626,N5633,N5640,N5647,N5654,N5718 
	,N5720,N5956,N5972,N5974,N5998,N6000,N6007,N6014 
	,N6021,N6028,N6035,N6042,N6049,N6056,N6063,N6070 
	,N6077,N6084,N6091,N6098,N6105,N6112,N6119,N6126 
	,N6133,N6140,N6147,N6154,N6299,N6304,N6430,N6439 
	,N6448,N6457,N6466,N6475,N6484,N6493,N6502,N6511 
	,N6520,N6529,N6538,N6547,N6565,N6574,N6583,N6592 
	,N6601,N6655,N6671,N6673,N6837,N6842,N6946,N7014 
	,N7038,N7040,N7068,N7070,N7083,N7091,N7099,N7128 
	,N7139,N7141,N7149,N7151,N7158,N7167,N7169,N7185 
	,N7187,N7203,N7205,N7221,N7223,N7230,N7239,N7241 
	,N7248,N7257,N7259,N7270,N7272,N7427,N7429,N7501 
	,N7505,N7661,N7663,N7931,N7933,N8017,N8100,N8102 
	,N8104,N8110,N8203,N8480,N8521,N8528,N8536,N8578 
	,N8941,N8990,N9246,N9251,N9260,N9267,N9274,N9281 
	,N9288,N9295,N9302,N9310,N9318,N9326,N9334,N9342 
	,N9350,N9358,N9366,N9374,N9382,N9390,N9398,N9404 
	,N9406,N9422,N9431,N9433,N9437,N9445,N9453,N9461 
	,N9469,N9477,N9485,N9493,N9501,N9509,N9517,N9525 
	,N9533,N9541,N9549,N9557,N9565,N9576,N10111,N10116 
	,N10123,N10157,N10159,N10166,N10168,N10173,N10175,N10193 
	,N10610,N10611,N10666,N10671;
reg x_reg_L1_12__retimed_I5171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5171_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23];
	end
assign N10193 = x_reg_L1_12__retimed_I5171_QOUT;
reg x_reg_L1_14__retimed_I5162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5162_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14];
	end
assign N10175 = x_reg_L1_14__retimed_I5162_QOUT;
reg x_reg_L1_20__retimed_I5161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5161_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20];
	end
assign N10173 = x_reg_L1_20__retimed_I5161_QOUT;
reg x_reg_L0_22__retimed_I5159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5159_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627;
	end
assign N10168 = x_reg_L0_22__retimed_I5159_QOUT;
reg x_reg_L0_22__retimed_I5158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5158_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596;
	end
assign N10166 = x_reg_L0_22__retimed_I5158_QOUT;
reg x_reg_L0_22__retimed_I5156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5156_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684;
	end
assign N10159 = x_reg_L0_22__retimed_I5156_QOUT;
reg x_reg_L0_22__retimed_I5155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5155_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706;
	end
assign N10157 = x_reg_L0_22__retimed_I5155_QOUT;
reg x_reg_L0_22__retimed_I5141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5141_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3];
	end
assign N10123 = x_reg_L0_22__retimed_I5141_QOUT;
reg x_reg_L0_22__retimed_I5139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5139_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
	end
assign N10116 = x_reg_L0_22__retimed_I5139_QOUT;
reg x_reg_L0_22__retimed_I5137_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5137_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4];
	end
assign N10111 = x_reg_L0_22__retimed_I5137_QOUT;
reg x_reg_L0_22__retimed_I4892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4892_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621;
	end
assign N9576 = x_reg_L0_22__retimed_I4892_QOUT;
reg x_reg_L0_22__retimed_I4888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4888_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719;
	end
assign N9565 = x_reg_L0_22__retimed_I4888_QOUT;
reg x_reg_L0_22__retimed_I4885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4885_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647;
	end
assign N9557 = x_reg_L0_22__retimed_I4885_QOUT;
reg x_reg_L0_22__retimed_I4882_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4882_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579;
	end
assign N9549 = x_reg_L0_22__retimed_I4882_QOUT;
reg x_reg_L0_22__retimed_I4879_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4879_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653;
	end
assign N9541 = x_reg_L0_22__retimed_I4879_QOUT;
reg x_reg_L0_22__retimed_I4876_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4876_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589;
	end
assign N9533 = x_reg_L0_22__retimed_I4876_QOUT;
reg x_reg_L0_22__retimed_I4873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4873_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663;
	end
assign N9525 = x_reg_L0_22__retimed_I4873_QOUT;
reg x_reg_L0_22__retimed_I4870_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4870_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595;
	end
assign N9517 = x_reg_L0_22__retimed_I4870_QOUT;
reg x_reg_L0_22__retimed_I4867_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4867_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673;
	end
assign N9509 = x_reg_L0_22__retimed_I4867_QOUT;
reg x_reg_L0_22__retimed_I4864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4864_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603;
	end
assign N9501 = x_reg_L0_22__retimed_I4864_QOUT;
reg x_reg_L0_22__retimed_I4861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4861_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679;
	end
assign N9493 = x_reg_L0_22__retimed_I4861_QOUT;
reg x_reg_L0_22__retimed_I4858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4858_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609;
	end
assign N9485 = x_reg_L0_22__retimed_I4858_QOUT;
reg x_reg_L0_22__retimed_I4855_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4855_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687;
	end
assign N9477 = x_reg_L0_22__retimed_I4855_QOUT;
reg x_reg_L0_22__retimed_I4852_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4852_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618;
	end
assign N9469 = x_reg_L0_22__retimed_I4852_QOUT;
reg x_reg_L0_22__retimed_I4849_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4849_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695;
	end
assign N9461 = x_reg_L0_22__retimed_I4849_QOUT;
reg x_reg_L0_22__retimed_I4846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4846_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626;
	end
assign N9453 = x_reg_L0_22__retimed_I4846_QOUT;
reg x_reg_L0_22__retimed_I4843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4843_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704;
	end
assign N9445 = x_reg_L0_22__retimed_I4843_QOUT;
reg x_reg_L0_22__retimed_I4840_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4840_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257;
	end
assign N9437 = x_reg_L0_22__retimed_I4840_QOUT;
reg x_reg_L0_22__retimed_I4839_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4839_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
	end
assign N9433 = x_reg_L0_22__retimed_I4839_QOUT;
reg x_reg_L0_22__retimed_I4838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4838_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613;
	end
assign N9431 = x_reg_L0_22__retimed_I4838_QOUT;
reg x_reg_L0_22__retimed_I4834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4834_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604;
	end
assign N9422 = x_reg_L0_22__retimed_I4834_QOUT;
reg x_reg_L0_22__retimed_I4829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4829_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604;
	end
assign N9406 = x_reg_L0_22__retimed_I4829_QOUT;
reg x_reg_L0_22__retimed_I4828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4828_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667;
	end
assign N9404 = x_reg_L0_22__retimed_I4828_QOUT;
reg x_reg_L0_22__retimed_I4827_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4827_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586;
	end
assign N9398 = x_reg_L0_22__retimed_I4827_QOUT;
reg x_reg_L0_22__retimed_I4825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4825_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668;
	end
assign N9390 = x_reg_L0_22__retimed_I4825_QOUT;
reg x_reg_L0_22__retimed_I4823_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4823_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648;
	end
assign N9382 = x_reg_L0_22__retimed_I4823_QOUT;
reg x_reg_L0_22__retimed_I4821_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4821_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713;
	end
assign N9374 = x_reg_L0_22__retimed_I4821_QOUT;
reg x_reg_L0_22__retimed_I4819_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4819_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628;
	end
assign N9366 = x_reg_L0_22__retimed_I4819_QOUT;
reg x_reg_L0_22__retimed_I4817_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4817_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692;
	end
assign N9358 = x_reg_L0_22__retimed_I4817_QOUT;
reg x_reg_L0_22__retimed_I4815_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4815_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610;
	end
assign N9350 = x_reg_L0_22__retimed_I4815_QOUT;
reg x_reg_L0_22__retimed_I4813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4813_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676;
	end
assign N9342 = x_reg_L0_22__retimed_I4813_QOUT;
reg x_reg_L0_22__retimed_I4811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4811_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593;
	end
assign N9334 = x_reg_L0_22__retimed_I4811_QOUT;
reg x_reg_L0_22__retimed_I4809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4809_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654;
	end
assign N9326 = x_reg_L0_22__retimed_I4809_QOUT;
reg x_reg_L0_22__retimed_I4807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4807_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722;
	end
assign N9318 = x_reg_L0_22__retimed_I4807_QOUT;
reg x_reg_L0_22__retimed_I4805_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4805_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636;
	end
assign N9310 = x_reg_L0_22__retimed_I4805_QOUT;
reg x_reg_L0_22__retimed_I4803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4803_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700;
	end
assign N9302 = x_reg_L0_22__retimed_I4803_QOUT;
reg x_reg_L0_22__retimed_I4801_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4801_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620;
	end
assign N9295 = x_reg_L0_22__retimed_I4801_QOUT;
reg x_reg_L0_22__retimed_I4799_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4799_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682;
	end
assign N9288 = x_reg_L0_22__retimed_I4799_QOUT;
reg x_reg_L0_22__retimed_I4797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4797_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600;
	end
assign N9281 = x_reg_L0_22__retimed_I4797_QOUT;
reg x_reg_L0_22__retimed_I4795_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4795_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665;
	end
assign N9274 = x_reg_L0_22__retimed_I4795_QOUT;
reg x_reg_L0_22__retimed_I4793_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4793_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582;
	end
assign N9267 = x_reg_L0_22__retimed_I4793_QOUT;
reg x_reg_L0_22__retimed_I4791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4791_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644;
	end
assign N9260 = x_reg_L0_22__retimed_I4791_QOUT;
reg x_reg_L0_22__retimed_I4788_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4788_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
	end
assign N9251 = x_reg_L0_22__retimed_I4788_QOUT;
reg x_reg_L0_22__retimed_I4787_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4787_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677;
	end
assign N9246 = x_reg_L0_22__retimed_I4787_QOUT;
reg x_reg_L0_22__retimed_I4696_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4696_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848;
	end
assign N8990 = x_reg_L0_22__retimed_I4696_QOUT;
reg x_reg_L0_22__retimed_I4678_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4678_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827;
	end
assign N8941 = x_reg_L0_22__retimed_I4678_QOUT;
reg x_reg_L0_22__retimed_I4607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4607_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486;
	end
assign N8578 = x_reg_L0_22__retimed_I4607_QOUT;
reg x_reg_L0_22__retimed_I4593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4593_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N8536 = x_reg_L0_22__retimed_I4593_QOUT;
reg x_reg_L0_22__retimed_I4590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4590_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N8528 = x_reg_L0_22__retimed_I4590_QOUT;
reg x_reg_L0_22__retimed_I4587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4587_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N8521 = x_reg_L0_22__retimed_I4587_QOUT;
reg x_reg_L0_22__retimed_I4570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4570_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N8480 = x_reg_L0_22__retimed_I4570_QOUT;
reg x_reg_L0_22__retimed_I4480_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4480_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N8203 = x_reg_L0_22__retimed_I4480_QOUT;
reg x_reg_L0_22__retimed_I4443_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4443_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N8110 = x_reg_L0_22__retimed_I4443_QOUT;
reg x_reg_L0_22__retimed_I4441_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4441_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N8104 = x_reg_L0_22__retimed_I4441_QOUT;
reg x_reg_L0_22__retimed_I4440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4440_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N8102 = x_reg_L0_22__retimed_I4440_QOUT;
reg x_reg_L0_22__retimed_I4439_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4439_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N8100 = x_reg_L0_22__retimed_I4439_QOUT;
reg x_reg_L0_22__retimed_I4406_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4406_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N8017 = x_reg_L0_22__retimed_I4406_QOUT;
reg x_reg_L1_21__retimed_I4373_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I4373_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23];
	end
assign N7933 = x_reg_L1_21__retimed_I4373_QOUT;
reg x_reg_L1_21__retimed_I4372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I4372_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564;
	end
assign N7931 = x_reg_L1_21__retimed_I4372_QOUT;
reg x_reg_L1_22__retimed_I4270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4270_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24];
	end
assign N7663 = x_reg_L1_22__retimed_I4270_QOUT;
reg x_reg_L1_22__retimed_I4269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I4269_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575;
	end
assign N7661 = x_reg_L1_22__retimed_I4269_QOUT;
reg x_reg_L1_12__retimed_I4208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4208_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
	end
assign N7505 = x_reg_L1_12__retimed_I4208_QOUT;
reg x_reg_L1_12__retimed_I4206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4206_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24];
	end
assign N7501 = x_reg_L1_12__retimed_I4206_QOUT;
reg x_reg_L1_12__retimed_I4178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4178_QOUT <= N7070;
	end
assign N7429 = x_reg_L1_12__retimed_I4178_QOUT;
reg x_reg_L1_12__retimed_I4177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4177_QOUT <= N7068;
	end
assign N7427 = x_reg_L1_12__retimed_I4177_QOUT;
reg x_reg_L1_23__retimed_I4115_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I4115_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
	end
assign N7272 = x_reg_L1_23__retimed_I4115_QOUT;
reg x_reg_L1_23__retimed_I4114_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I4114_QOUT <= N7248;
	end
assign N7270 = x_reg_L1_23__retimed_I4114_QOUT;
reg x_reg_L1_24__retimed_I4111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I4111_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135;
	end
assign N7259 = x_reg_L1_24__retimed_I4111_QOUT;
reg x_reg_L1_24__retimed_I4110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I4110_QOUT <= N7230;
	end
assign N7257 = x_reg_L1_24__retimed_I4110_QOUT;
reg x_reg_L0_22__retimed_I4107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4107_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N7248 = x_reg_L0_22__retimed_I4107_QOUT;
reg x_reg_L1_25__retimed_I4105_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I4105_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
	end
assign N7241 = x_reg_L1_25__retimed_I4105_QOUT;
reg x_reg_L1_25__retimed_I4104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I4104_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729;
	end
assign N7239 = x_reg_L1_25__retimed_I4104_QOUT;
reg x_reg_L0_22__retimed_I4101_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4101_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738;
	end
assign N7230 = x_reg_L0_22__retimed_I4101_QOUT;
reg x_reg_L1_26__retimed_I4099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I4099_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754;
	end
assign N7223 = x_reg_L1_26__retimed_I4099_QOUT;
reg x_reg_L1_26__retimed_I4098_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I4098_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270;
	end
assign N7221 = x_reg_L1_26__retimed_I4098_QOUT;
reg x_reg_L1_27__retimed_I4093_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I4093_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142;
	end
assign N7205 = x_reg_L1_27__retimed_I4093_QOUT;
reg x_reg_L1_27__retimed_I4092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I4092_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724;
	end
assign N7203 = x_reg_L1_27__retimed_I4092_QOUT;
reg x_reg_L1_28__retimed_I4087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I4087_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736;
	end
assign N7187 = x_reg_L1_28__retimed_I4087_QOUT;
reg x_reg_L1_28__retimed_I4086_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I4086_QOUT <= N7158;
	end
assign N7185 = x_reg_L1_28__retimed_I4086_QOUT;
reg x_reg_L1_29__retimed_I4081_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I4081_QOUT <= N7141;
	end
assign N7169 = x_reg_L1_29__retimed_I4081_QOUT;
reg x_reg_L1_29__retimed_I4080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I4080_QOUT <= N7139;
	end
assign N7167 = x_reg_L1_29__retimed_I4080_QOUT;
reg x_reg_L0_22__retimed_I4077_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4077_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
	end
assign N7158 = x_reg_L0_22__retimed_I4077_QOUT;
reg x_reg_L1_30__retimed_I4075_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I4075_QOUT <= N7128;
	end
assign N7151 = x_reg_L1_30__retimed_I4075_QOUT;
reg x_reg_L1_30__retimed_I4074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I4074_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446;
	end
assign N7149 = x_reg_L1_30__retimed_I4074_QOUT;
reg x_reg_L0_22__retimed_I4072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4072_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439;
	end
assign N7141 = x_reg_L0_22__retimed_I4072_QOUT;
reg x_reg_L0_22__retimed_I4071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N7139 = x_reg_L0_22__retimed_I4071_QOUT;
reg x_reg_L0_22__retimed_I4068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N7128 = x_reg_L0_22__retimed_I4068_QOUT;
reg x_reg_L1_12__retimed_I4058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4058_QOUT <= N7014;
	end
assign N7099 = x_reg_L1_12__retimed_I4058_QOUT;
reg x_reg_L1_12__retimed_I4056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4056_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742;
	end
assign N7091 = x_reg_L1_12__retimed_I4056_QOUT;
reg x_reg_L1_12__retimed_I4053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4053_QOUT <= N10116;
	end
assign N7083 = x_reg_L1_12__retimed_I4053_QOUT;
reg x_reg_L0_22__retimed_I4049_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4049_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2];
	end
assign N7070 = x_reg_L0_22__retimed_I4049_QOUT;
reg x_reg_L0_22__retimed_I4048_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4048_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N7068 = x_reg_L0_22__retimed_I4048_QOUT;
reg x_reg_L1_12__retimed_I4036_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4036_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5];
	end
assign N7040 = x_reg_L1_12__retimed_I4036_QOUT;
reg x_reg_L1_12__retimed_I4035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I4035_QOUT <= N6946;
	end
assign N7038 = x_reg_L1_12__retimed_I4035_QOUT;
reg x_reg_L0_22__retimed_I4026_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I4026_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707;
	end
assign N7014 = x_reg_L0_22__retimed_I4026_QOUT;
reg x_reg_L0_22__retimed_I3999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3999_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681;
	end
assign N6946 = x_reg_L0_22__retimed_I3999_QOUT;
reg x_reg_L1_23__retimed_I3965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3965_QOUT <= N6304;
	end
assign N6842 = x_reg_L1_23__retimed_I3965_QOUT;
reg x_reg_L1_22__retimed_I3963_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3963_QOUT <= N6299;
	end
assign N6837 = x_reg_L1_22__retimed_I3963_QOUT;
reg x_reg_L1_23__retimed_I3927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3927_QOUT <= N5974;
	end
assign N6673 = x_reg_L1_23__retimed_I3927_QOUT;
reg x_reg_L1_23__retimed_I3926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I3926_QOUT <= N5972;
	end
assign N6671 = x_reg_L1_23__retimed_I3926_QOUT;
reg x_reg_L1_22__retimed_I3923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I3923_QOUT <= N5956;
	end
assign N6655 = x_reg_L1_22__retimed_I3923_QOUT;
reg x_reg_L1_19__retimed_I3909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3909_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19];
	end
assign N6601 = x_reg_L1_19__retimed_I3909_QOUT;
reg x_reg_L1_18__retimed_I3905_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3905_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18];
	end
assign N6592 = x_reg_L1_18__retimed_I3905_QOUT;
reg x_reg_L1_17__retimed_I3901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3901_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17];
	end
assign N6583 = x_reg_L1_17__retimed_I3901_QOUT;
reg x_reg_L1_16__retimed_I3897_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3897_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16];
	end
assign N6574 = x_reg_L1_16__retimed_I3897_QOUT;
reg x_reg_L1_15__retimed_I3893_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3893_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15];
	end
assign N6565 = x_reg_L1_15__retimed_I3893_QOUT;
reg x_reg_L1_13__retimed_I3885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3885_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13];
	end
assign N6547 = x_reg_L1_13__retimed_I3885_QOUT;
reg x_reg_L1_12__retimed_I3881_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3881_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12];
	end
assign N6538 = x_reg_L1_12__retimed_I3881_QOUT;
reg x_reg_L1_11__retimed_I3877_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3877_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11];
	end
assign N6529 = x_reg_L1_11__retimed_I3877_QOUT;
reg x_reg_L1_10__retimed_I3873_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3873_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10];
	end
assign N6520 = x_reg_L1_10__retimed_I3873_QOUT;
reg x_reg_L1_9__retimed_I3869_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3869_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9];
	end
assign N6511 = x_reg_L1_9__retimed_I3869_QOUT;
reg x_reg_L1_8__retimed_I3865_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3865_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8];
	end
assign N6502 = x_reg_L1_8__retimed_I3865_QOUT;
reg x_reg_L1_7__retimed_I3861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3861_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7];
	end
assign N6493 = x_reg_L1_7__retimed_I3861_QOUT;
reg x_reg_L1_6__retimed_I3857_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3857_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6];
	end
assign N6484 = x_reg_L1_6__retimed_I3857_QOUT;
reg x_reg_L1_5__retimed_I3853_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3853_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5];
	end
assign N6475 = x_reg_L1_5__retimed_I3853_QOUT;
reg x_reg_L1_4__retimed_I3849_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3849_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4];
	end
assign N6466 = x_reg_L1_4__retimed_I3849_QOUT;
reg x_reg_L1_3__retimed_I3845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3845_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3];
	end
assign N6457 = x_reg_L1_3__retimed_I3845_QOUT;
reg x_reg_L1_2__retimed_I3841_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3841_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2];
	end
assign N6448 = x_reg_L1_2__retimed_I3841_QOUT;
reg x_reg_L1_1__retimed_I3837_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3837_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1];
	end
assign N6439 = x_reg_L1_1__retimed_I3837_QOUT;
reg x_reg_L1_0__retimed_I3833_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3833_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0];
	end
assign N6430 = x_reg_L1_0__retimed_I3833_QOUT;
reg x_reg_L0_23__retimed_I3782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3782_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N6304 = x_reg_L0_23__retimed_I3782_QOUT;
reg x_reg_L0_7__retimed_I3780_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3780_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912;
	end
assign N6299 = x_reg_L0_7__retimed_I3780_QOUT;
reg x_reg_L1_0__retimed_I3747_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I3747_QOUT <= N5654;
	end
assign N6154 = x_reg_L1_0__retimed_I3747_QOUT;
reg x_reg_L1_1__retimed_I3744_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I3744_QOUT <= N5647;
	end
assign N6147 = x_reg_L1_1__retimed_I3744_QOUT;
reg x_reg_L1_2__retimed_I3741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I3741_QOUT <= N5640;
	end
assign N6140 = x_reg_L1_2__retimed_I3741_QOUT;
reg x_reg_L1_3__retimed_I3738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I3738_QOUT <= N5633;
	end
assign N6133 = x_reg_L1_3__retimed_I3738_QOUT;
reg x_reg_L1_4__retimed_I3735_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I3735_QOUT <= N5626;
	end
assign N6126 = x_reg_L1_4__retimed_I3735_QOUT;
reg x_reg_L1_5__retimed_I3732_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I3732_QOUT <= N5619;
	end
assign N6119 = x_reg_L1_5__retimed_I3732_QOUT;
reg x_reg_L1_6__retimed_I3729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I3729_QOUT <= N5612;
	end
assign N6112 = x_reg_L1_6__retimed_I3729_QOUT;
reg x_reg_L1_7__retimed_I3726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I3726_QOUT <= N5605;
	end
assign N6105 = x_reg_L1_7__retimed_I3726_QOUT;
reg x_reg_L1_8__retimed_I3723_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I3723_QOUT <= N5598;
	end
assign N6098 = x_reg_L1_8__retimed_I3723_QOUT;
reg x_reg_L1_9__retimed_I3720_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I3720_QOUT <= N5591;
	end
assign N6091 = x_reg_L1_9__retimed_I3720_QOUT;
reg x_reg_L1_10__retimed_I3717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I3717_QOUT <= N5584;
	end
assign N6084 = x_reg_L1_10__retimed_I3717_QOUT;
reg x_reg_L1_11__retimed_I3714_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I3714_QOUT <= N5577;
	end
assign N6077 = x_reg_L1_11__retimed_I3714_QOUT;
reg x_reg_L1_12__retimed_I3711_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I3711_QOUT <= N5570;
	end
assign N6070 = x_reg_L1_12__retimed_I3711_QOUT;
reg x_reg_L1_13__retimed_I3708_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I3708_QOUT <= N5563;
	end
assign N6063 = x_reg_L1_13__retimed_I3708_QOUT;
reg x_reg_L1_14__retimed_I3705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I3705_QOUT <= N5556;
	end
assign N6056 = x_reg_L1_14__retimed_I3705_QOUT;
reg x_reg_L1_15__retimed_I3702_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I3702_QOUT <= N5549;
	end
assign N6049 = x_reg_L1_15__retimed_I3702_QOUT;
reg x_reg_L1_16__retimed_I3699_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I3699_QOUT <= N5542;
	end
assign N6042 = x_reg_L1_16__retimed_I3699_QOUT;
reg x_reg_L1_17__retimed_I3696_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I3696_QOUT <= N5535;
	end
assign N6035 = x_reg_L1_17__retimed_I3696_QOUT;
reg x_reg_L1_18__retimed_I3693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I3693_QOUT <= N5528;
	end
assign N6028 = x_reg_L1_18__retimed_I3693_QOUT;
reg x_reg_L1_19__retimed_I3690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I3690_QOUT <= N5521;
	end
assign N6021 = x_reg_L1_19__retimed_I3690_QOUT;
reg x_reg_L1_20__retimed_I3687_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I3687_QOUT <= N5514;
	end
assign N6014 = x_reg_L1_20__retimed_I3687_QOUT;
reg x_reg_L1_21__retimed_I3684_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I3684_QOUT <= N5507;
	end
assign N6007 = x_reg_L1_21__retimed_I3684_QOUT;
reg x_reg_L0_31__retimed_I3681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3681_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N6000 = x_reg_L0_31__retimed_I3681_QOUT;
reg x_reg_L0_31__retimed_I3680_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3680_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5998 = x_reg_L0_31__retimed_I3680_QOUT;
reg x_reg_L0_23__retimed_I3672_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3672_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5974 = x_reg_L0_23__retimed_I3672_QOUT;
reg x_reg_L0_23__retimed_I3671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I3671_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5972 = x_reg_L0_23__retimed_I3671_QOUT;
reg x_reg_L0_22__retimed_I3668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I3668_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5956 = x_reg_L0_22__retimed_I3668_QOUT;
reg x_reg_L0_31__retimed_I3573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3573_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113;
	end
assign N5720 = x_reg_L0_31__retimed_I3573_QOUT;
reg x_reg_L0_31__retimed_I3572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__retimed_I3572_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122;
	end
assign N5718 = x_reg_L0_31__retimed_I3572_QOUT;
reg x_reg_L0_0__retimed_I3545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I3545_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5654 = x_reg_L0_0__retimed_I3545_QOUT;
reg x_reg_L0_1__retimed_I3542_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I3542_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5647 = x_reg_L0_1__retimed_I3542_QOUT;
reg x_reg_L0_2__retimed_I3539_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I3539_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5640 = x_reg_L0_2__retimed_I3539_QOUT;
reg x_reg_L0_3__retimed_I3536_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I3536_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5633 = x_reg_L0_3__retimed_I3536_QOUT;
reg x_reg_L0_4__retimed_I3533_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I3533_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5626 = x_reg_L0_4__retimed_I3533_QOUT;
reg x_reg_L0_5__retimed_I3530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I3530_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5619 = x_reg_L0_5__retimed_I3530_QOUT;
reg x_reg_L0_6__retimed_I3527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I3527_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5612 = x_reg_L0_6__retimed_I3527_QOUT;
reg x_reg_L0_7__retimed_I3524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I3524_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5605 = x_reg_L0_7__retimed_I3524_QOUT;
reg x_reg_L0_8__retimed_I3521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I3521_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5598 = x_reg_L0_8__retimed_I3521_QOUT;
reg x_reg_L0_9__retimed_I3518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I3518_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5591 = x_reg_L0_9__retimed_I3518_QOUT;
reg x_reg_L0_10__retimed_I3515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I3515_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5584 = x_reg_L0_10__retimed_I3515_QOUT;
reg x_reg_L0_11__retimed_I3512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I3512_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5577 = x_reg_L0_11__retimed_I3512_QOUT;
reg x_reg_L0_12__retimed_I3509_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I3509_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5570 = x_reg_L0_12__retimed_I3509_QOUT;
reg x_reg_L0_13__retimed_I3506_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I3506_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5563 = x_reg_L0_13__retimed_I3506_QOUT;
reg x_reg_L0_14__retimed_I3503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I3503_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5556 = x_reg_L0_14__retimed_I3503_QOUT;
reg x_reg_L0_15__retimed_I3500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I3500_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5549 = x_reg_L0_15__retimed_I3500_QOUT;
reg x_reg_L0_16__retimed_I3497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I3497_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5542 = x_reg_L0_16__retimed_I3497_QOUT;
reg x_reg_L0_17__retimed_I3494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I3494_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5535 = x_reg_L0_17__retimed_I3494_QOUT;
reg x_reg_L0_18__retimed_I3491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I3491_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5528 = x_reg_L0_18__retimed_I3491_QOUT;
reg x_reg_L0_19__retimed_I3488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I3488_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5521 = x_reg_L0_19__retimed_I3488_QOUT;
reg x_reg_L0_20__retimed_I3485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I3485_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5514 = x_reg_L0_20__retimed_I3485_QOUT;
reg x_reg_L0_21__retimed_I3482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I3482_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5507 = x_reg_L0_21__retimed_I3482_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123 = !(((a_man[0] | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168 = !(b_exp[0] & b_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202 = !((b_exp[7] & b_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056 = !(a_exp[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544 = !a_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426 = !(b_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479 = !(b_man[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410 = !a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530 = !(b_man[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433 = !(b_man[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485 = !(b_man[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537 = !(b_man[16] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489 = !a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496 = !(b_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550 = !(b_man[10] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451 = !(b_man[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453 = !a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439 = !(b_man[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492 = !(b_man[14] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542 = !(b_man[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446 = !(b_man[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503 = !(b_man[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525 = !a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404 = !(b_man[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455 = !(b_man[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547 = !a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506 = !(b_man[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408 = !(b_man[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460 = !(b_man[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449 = !(b_man[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527 = !(((a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546 = !(b_man[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494 = !(b_man[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443 = !(b_man[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540 = !(b_man[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488 = !(b_man[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437 = !(b_man[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534 = !(b_man[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483 = !(b_man[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430 = !(b_man[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528 = !(b_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477 = !(b_man[12] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424 = !(b_man[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524 = !(b_man[14] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471 = !(b_man[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419 = !(b_man[16] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518 = !(b_man[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465 = !(b_man[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413 = !(b_man[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511 = !(b_man[20] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459 = !(b_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475) | (b_man[22] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565} = {1'B0, a_exp[0]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563} + {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556 ^ a_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[11]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[13]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[4]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[4]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149) & a_man[3]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769 & a_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353)) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150) & a_man[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635 = !(N10166 | N10168);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635 | (!N9398));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606 = !(N9576 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718 = (!N9565) | (N9382 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709 = (!N9557) | (N9374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709) ^ N9366;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718) ^ N9374;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643) ^ N9382;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611 = !N10168;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611) | (N9431 & N9433);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635) ^ N9398;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864);
assign N10666 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667 = !N10666;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691 = (!N9422) | (N9406 & N9404);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691) ^ N9390;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!N9404) ^ N9406;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] = (!N10157) ^ N10159;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | N8521);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[13]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[12]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148) & a_man[9]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612 = (!N9549) | (N9366 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583 = (!N9541) | (N9358 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616 = (!N9533) | (N9350 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717 = (!N9525) | (N9342 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585 = (!N9517) | (N9334 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664 = (!N9509) | (N9326 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659 = (!N9501) | (N9318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723 = (!N9493) | (N9310 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723) ^ N9302;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659) ^ N9310;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664) ^ N9318;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585) ^ N9326;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717) ^ N9334;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616) ^ N9342;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583) ^ N9350;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612) ^ N9358;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147) & a_man[17]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699 = (!N9485) | (N9302 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597 = (!N9477) | (N9295 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701 = (!N9469) | (N9288 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578 = (!N9461) | (N9281 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578) ^ N9274;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701) ^ N9281;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597) ^ N9288;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699) ^ N9295;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666 = (!N9453) | (N9274 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672 = (!N9445) | (N9267 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672) ^ N9260;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666) ^ N9267;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594 = (!N9437) | (N9260 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624 = !(N9246 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] = N9251 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594) ^ N9246;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[2]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729} = {1'B0, N7068} + {1'B0, N7070};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3] | (!N8521));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863 = !((N8990 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4860) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4881);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4902);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4889) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4911);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4824)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4838)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4866);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4877) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4917);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0] = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 = !(N8941 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831 & (!N8941));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4828;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285 = N8521 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214 = N8528 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143 = N8536 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5284 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179) & N8536);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5269 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N8521);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5233 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178) & N8528);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8182 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32 & a_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32) & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631 = N8578 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N8480) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280 = !(N8017 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & N8110) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633 = N8203 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269 = !(((N8100 | N8102) | N8104) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5576 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8080;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8086;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8139;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]} = {1'B0, N7270} + {1'B0, N7272} + {1'B0, N10193};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]} = {1'B0, N7257} + {1'B0, N7259} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13744};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]} = {1'B0, N7239} + {1'B0, N7241} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13695};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[3]);
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754} = {1'B0, N10123} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724} = {1'B0, N10111} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]} = {1'B0, N7221} + {1'B0, N7223} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13732};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]} = {1'B0, N7203} + {1'B0, N7205} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13685};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]} = {1'B0, N7185} + {1'B0, N7187} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13722};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 & a_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433) & b_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]} = {1'B0, N7167} + {1'B0, N7169} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13746};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433 & a_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433) & b_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742 = !N10116;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446 = !N10116;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686} = {1'B0, N7149} + {1'B0, N7151} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734;
assign N10610 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710;
assign N10611 = !N10610;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683 = !(N7091 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730 = !(N7091 & N10611);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13699 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13738) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13730);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642 = (N10193 & N7501) | N7505;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754 = !((N7427 & N7429) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62 = !(N7099 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740 = !(N7083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701 = !(((N7038 | N7040) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13740);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13692 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13719) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13706) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13701);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__71;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 | (!N6655));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70 = N6837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 = !(N6655 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22] = (!N7661) ^ N7663;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21] = N7931 ^ N7933;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6007);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & N10173));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6014);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & N6601));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6021);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184 & N6592));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6028);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & N6583));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6035);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & N6574));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6042);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & N6565));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6049);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & N10175));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6056);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185 & N6547));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6063);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & N6538));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6070);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & N6529));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6077);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & N6520));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6084);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & N6511));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6091);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186 & N6502));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6098);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6493));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6105);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594 = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6484));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6112);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6475));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6466));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6126);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6457));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6133);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3] & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6448));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6140);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6439));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6147);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_man[0]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2] ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188 & N6430));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942 & N6154);
assign N10671 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7] = !N10671;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869 = ((N6673 | N6671) | N6655) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651 = N6842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0] = ((N6671 | N6673) | N6655) | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5] & N6000) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]) & N5998);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31] = (N5718 & fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116) | ((!N5718) & N5720);
reg x_reg_L1_31__I1159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1159_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_L1_31__I1159_QOUT;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLjwTADZrRo= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



