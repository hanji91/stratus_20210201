/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:09 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794,
	float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796;
wire N5603,N5608,N5613,N5618,N5623,N5628,N5633 
	,N5638,N5643,N11736,N11738,N11899,N11904,N11909,N11914 
	,N11919,N11924,N11929,N12012,N12014,N12065,N12067,N12072 
	,N12077,N12082,N12087,N12092,N12095,N12097,N12110,N12112 
	,N12118,N12120,N12136,N12138,N12144,N12146,N12154,N12156 
	,N12166,N12168,N12176,N12178,N12184,N12186,N12194,N12196 
	,N12206,N12268,N12270,N12272,N12294,N12298,N12320,N12354 
	,N12356,N12386,N12388,N12418,N12450,N12460,N12464,N12466 
	,N12538,N12586,N12599,N12605,N12607,N12609,N12647,N12669 
	,N12671,N12673,N12731,N12744,N12746,N12748,N12753,N12807 
	,N12823,N12825,N12827,N12885,N12893,N12895,N12897,N12963 
	,N13000,N13002,N13004,N13074,N13081,N13087,N13089,N13091 
	,N13094,N13104,N13189,N13197,N13199,N13201,N13205,N13207 
	,N13209,N13218,N13220,N13222,N13225,N13227,N13305,N13311 
	,N13319,N13335,N13337,N13424,N13430,N13432,N13436,N13448 
	,N13458,N13460,N13462,N13466,N13500,N13523,N13541,N13549 
	,N13551,N13555,N13557,N13583,N13585,N13587,N13591,N13593 
	,N13599,N13601,N13607,N13609,N13611,N13630,N13647,N13649 
	,N13659,N13673,N13675,N13681,N13685,N13689,N13693,N13697 
	,N13699,N13709,N13712,N13718,N13720,N13722,N13725,N13731 
	,N13733,N13735,N13761,N13763,N13769,N13771,N13773,N13777 
	,N13779,N13785,N13787,N13789,N13798,N13800,N13802,N13806 
	,N13808,N13810,N13822,N13824,N13835,N13837,N13842,N13852 
	,N13854,N13856,N13862,N13864,N13866,N13870,N13872,N13874 
	,N13878,N13880,N13882,N13888,N13890,N13892,N13896,N13898 
	,N13900,N14500,N14505,N14510,N14513,N14518,N14523,N14528 
	,N14533;
reg x_reg_L0_22__retimed_I7921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7921_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355;
	end
assign N14533 = x_reg_L0_22__retimed_I7921_QOUT;
reg x_reg_L0_22__retimed_I7919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7919_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205;
	end
assign N14528 = x_reg_L0_22__retimed_I7919_QOUT;
reg x_reg_L0_22__retimed_I7917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7917_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132;
	end
assign N14523 = x_reg_L0_22__retimed_I7917_QOUT;
reg x_reg_L0_22__retimed_I7915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7915_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397;
	end
assign N14518 = x_reg_L0_22__retimed_I7915_QOUT;
reg x_reg_L0_22__retimed_I7913_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7913_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164;
	end
assign N14513 = x_reg_L0_22__retimed_I7913_QOUT;
reg x_reg_L0_22__retimed_I7912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7912_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219;
	end
assign N14510 = x_reg_L0_22__retimed_I7912_QOUT;
reg x_reg_L0_22__retimed_I7910_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7910_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365;
	end
assign N14505 = x_reg_L0_22__retimed_I7910_QOUT;
reg x_reg_L0_22__retimed_I7908_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7908_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292;
	end
assign N14500 = x_reg_L0_22__retimed_I7908_QOUT;
reg x_reg_L0_22__retimed_I7660_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7660_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[8];
	end
assign N13900 = x_reg_L0_22__retimed_I7660_QOUT;
reg x_reg_L0_22__retimed_I7659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7659_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[8];
	end
assign N13898 = x_reg_L0_22__retimed_I7659_QOUT;
reg x_reg_L0_22__retimed_I7658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7658_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[8];
	end
assign N13896 = x_reg_L0_22__retimed_I7658_QOUT;
reg x_reg_L0_22__retimed_I7657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7657_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949;
	end
assign N13892 = x_reg_L0_22__retimed_I7657_QOUT;
reg x_reg_L0_22__retimed_I7656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7656_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[7];
	end
assign N13890 = x_reg_L0_22__retimed_I7656_QOUT;
reg x_reg_L0_22__retimed_I7655_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7655_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445;
	end
assign N13888 = x_reg_L0_22__retimed_I7655_QOUT;
reg x_reg_L0_22__retimed_I7654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7654_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178;
	end
assign N13882 = x_reg_L0_22__retimed_I7654_QOUT;
reg x_reg_L0_22__retimed_I7653_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7653_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338;
	end
assign N13880 = x_reg_L0_22__retimed_I7653_QOUT;
reg x_reg_L0_22__retimed_I7652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7652_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371;
	end
assign N13878 = x_reg_L0_22__retimed_I7652_QOUT;
reg x_reg_L0_22__retimed_I7651_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7651_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075;
	end
assign N13874 = x_reg_L0_22__retimed_I7651_QOUT;
reg x_reg_L0_22__retimed_I7650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7650_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264;
	end
assign N13872 = x_reg_L0_22__retimed_I7650_QOUT;
reg x_reg_L0_22__retimed_I7649_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7649_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233;
	end
assign N13870 = x_reg_L0_22__retimed_I7649_QOUT;
reg x_reg_L0_22__retimed_I7648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7648_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[9];
	end
assign N13866 = x_reg_L0_22__retimed_I7648_QOUT;
reg x_reg_L0_22__retimed_I7647_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7647_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[9];
	end
assign N13864 = x_reg_L0_22__retimed_I7647_QOUT;
reg x_reg_L0_22__retimed_I7646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7646_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[9];
	end
assign N13862 = x_reg_L0_22__retimed_I7646_QOUT;
reg x_reg_L0_22__retimed_I7644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7644_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789;
	end
assign N13856 = x_reg_L0_22__retimed_I7644_QOUT;
reg x_reg_L0_22__retimed_I7643_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7643_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528;
	end
assign N13854 = x_reg_L0_22__retimed_I7643_QOUT;
reg x_reg_L0_22__retimed_I7642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7642_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623;
	end
assign N13852 = x_reg_L0_22__retimed_I7642_QOUT;
reg x_reg_L0_22__retimed_I7638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7638_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925;
	end
assign N13842 = x_reg_L0_22__retimed_I7638_QOUT;
reg x_reg_L0_22__retimed_I7636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7636_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839;
	end
assign N13837 = x_reg_L0_22__retimed_I7636_QOUT;
reg x_reg_L0_22__retimed_I7635_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7635_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[8];
	end
assign N13835 = x_reg_L0_22__retimed_I7635_QOUT;
reg x_reg_L0_22__retimed_I7632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7632_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588;
	end
assign N13824 = x_reg_L0_22__retimed_I7632_QOUT;
reg x_reg_L0_22__retimed_I7631_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7631_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802;
	end
assign N13822 = x_reg_L0_22__retimed_I7631_QOUT;
reg x_reg_L0_22__retimed_I7630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7630_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236;
	end
assign N13810 = x_reg_L0_22__retimed_I7630_QOUT;
reg x_reg_L0_22__retimed_I7629_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7629_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372;
	end
assign N13808 = x_reg_L0_22__retimed_I7629_QOUT;
reg x_reg_L0_22__retimed_I7628_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7628_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166;
	end
assign N13806 = x_reg_L0_22__retimed_I7628_QOUT;
reg x_reg_L0_22__retimed_I7627_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7627_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363;
	end
assign N13802 = x_reg_L0_22__retimed_I7627_QOUT;
reg x_reg_L0_22__retimed_I7626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7626_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158;
	end
assign N13800 = x_reg_L0_22__retimed_I7626_QOUT;
reg x_reg_L0_22__retimed_I7625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7625_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291;
	end
assign N13798 = x_reg_L0_22__retimed_I7625_QOUT;
reg x_reg_L0_22__retimed_I7622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7622_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378;
	end
assign N13789 = x_reg_L0_22__retimed_I7622_QOUT;
reg x_reg_L0_22__retimed_I7621_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7621_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304;
	end
assign N13787 = x_reg_L0_22__retimed_I7621_QOUT;
reg x_reg_L0_22__retimed_I7620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7620_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172;
	end
assign N13785 = x_reg_L0_22__retimed_I7620_QOUT;
reg x_reg_L0_22__retimed_I7618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7618_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[10];
	end
assign N13779 = x_reg_L0_22__retimed_I7618_QOUT;
reg x_reg_L0_22__retimed_I7617_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7617_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[10];
	end
assign N13777 = x_reg_L0_22__retimed_I7617_QOUT;
reg x_reg_L0_22__retimed_I7616_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7616_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388;
	end
assign N13773 = x_reg_L0_22__retimed_I7616_QOUT;
reg x_reg_L0_22__retimed_I7615_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7615_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238;
	end
assign N13771 = x_reg_L0_22__retimed_I7615_QOUT;
reg x_reg_L0_22__retimed_I7614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7614_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062;
	end
assign N13769 = x_reg_L0_22__retimed_I7614_QOUT;
reg x_reg_L0_22__retimed_I7612_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7612_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327;
	end
assign N13763 = x_reg_L0_22__retimed_I7612_QOUT;
reg x_reg_L0_22__retimed_I7611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7611_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151;
	end
assign N13761 = x_reg_L0_22__retimed_I7611_QOUT;
reg x_reg_L0_22__retimed_I7602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7602_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844;
	end
assign N13735 = x_reg_L0_22__retimed_I7602_QOUT;
reg x_reg_L0_22__retimed_I7601_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7601_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330;
	end
assign N13733 = x_reg_L0_22__retimed_I7601_QOUT;
reg x_reg_L0_22__retimed_I7600_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7600_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206;
	end
assign N13731 = x_reg_L0_22__retimed_I7600_QOUT;
reg x_reg_L0_22__retimed_I7598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7598_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322;
	end
assign N13725 = x_reg_L0_22__retimed_I7598_QOUT;
reg x_reg_L0_22__retimed_I7597_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7597_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112;
	end
assign N13722 = x_reg_L0_22__retimed_I7597_QOUT;
reg x_reg_L0_22__retimed_I7596_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7596_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123;
	end
assign N13720 = x_reg_L0_22__retimed_I7596_QOUT;
reg x_reg_L0_22__retimed_I7595_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7595_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313;
	end
assign N13718 = x_reg_L0_22__retimed_I7595_QOUT;
reg x_reg_L0_22__retimed_I7593_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7593_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246;
	end
assign N13712 = x_reg_L0_22__retimed_I7593_QOUT;
reg x_reg_L0_22__retimed_I7592_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7592_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179;
	end
assign N13709 = x_reg_L0_22__retimed_I7592_QOUT;
reg x_reg_L0_22__retimed_I7588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7588_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184;
	end
assign N13699 = x_reg_L0_22__retimed_I7588_QOUT;
reg x_reg_L0_22__retimed_I7587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7587_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320;
	end
assign N13697 = x_reg_L0_22__retimed_I7587_QOUT;
reg x_reg_L0_22__retimed_I7586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7586_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203;
	end
assign N13693 = x_reg_L0_22__retimed_I7586_QOUT;
reg x_reg_L0_22__retimed_I7584_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7584_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395;
	end
assign N13689 = x_reg_L0_22__retimed_I7584_QOUT;
reg x_reg_L0_22__retimed_I7583_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7583_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069;
	end
assign N13685 = x_reg_L0_22__retimed_I7583_QOUT;
reg x_reg_L0_22__retimed_I7581_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7581_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269;
	end
assign N13681 = x_reg_L0_22__retimed_I7581_QOUT;
reg x_reg_L0_22__retimed_I7579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7579_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144;
	end
assign N13675 = x_reg_L0_22__retimed_I7579_QOUT;
reg x_reg_L0_22__retimed_I7578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7578_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130;
	end
assign N13673 = x_reg_L0_22__retimed_I7578_QOUT;
reg x_reg_L0_22__retimed_I7573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7573_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150;
	end
assign N13659 = x_reg_L0_22__retimed_I7573_QOUT;
reg x_reg_L0_22__retimed_I7569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7569_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[11];
	end
assign N13649 = x_reg_L0_22__retimed_I7569_QOUT;
reg x_reg_L0_22__retimed_I7568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7568_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[11];
	end
assign N13647 = x_reg_L0_22__retimed_I7568_QOUT;
reg x_reg_L0_22__retimed_I7561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7561_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197;
	end
assign N13630 = x_reg_L0_22__retimed_I7561_QOUT;
reg x_reg_L0_22__retimed_I7555_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7555_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044;
	end
assign N13611 = x_reg_L0_22__retimed_I7555_QOUT;
reg x_reg_L0_22__retimed_I7554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7554_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030;
	end
assign N13609 = x_reg_L0_22__retimed_I7554_QOUT;
reg x_reg_L0_22__retimed_I7553_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7553_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535;
	end
assign N13607 = x_reg_L0_22__retimed_I7553_QOUT;
reg x_reg_L0_22__retimed_I7551_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7551_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198;
	end
assign N13601 = x_reg_L0_22__retimed_I7551_QOUT;
reg x_reg_L0_22__retimed_I7550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7550_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133;
	end
assign N13599 = x_reg_L0_22__retimed_I7550_QOUT;
reg x_reg_L0_22__retimed_I7548_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7548_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122;
	end
assign N13593 = x_reg_L0_22__retimed_I7548_QOUT;
reg x_reg_L0_22__retimed_I7547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7547_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389;
	end
assign N13591 = x_reg_L0_22__retimed_I7547_QOUT;
reg x_reg_L0_22__retimed_I7546_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7546_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762;
	end
assign N13587 = x_reg_L0_22__retimed_I7546_QOUT;
reg x_reg_L0_22__retimed_I7545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7545_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246;
	end
assign N13585 = x_reg_L0_22__retimed_I7545_QOUT;
reg x_reg_L0_22__retimed_I7544_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7544_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231;
	end
assign N13583 = x_reg_L0_22__retimed_I7544_QOUT;
reg x_reg_L0_22__retimed_I7534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7534_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396;
	end
assign N13557 = x_reg_L0_22__retimed_I7534_QOUT;
reg x_reg_L0_22__retimed_I7533_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7533_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260;
	end
assign N13555 = x_reg_L0_22__retimed_I7533_QOUT;
reg x_reg_L0_22__retimed_I7532_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7532_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370;
	end
assign N13551 = x_reg_L0_22__retimed_I7532_QOUT;
reg x_reg_L0_22__retimed_I7531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7531_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223;
	end
assign N13549 = x_reg_L0_22__retimed_I7531_QOUT;
reg x_reg_L0_22__retimed_I7528_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7528_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311;
	end
assign N13541 = x_reg_L0_22__retimed_I7528_QOUT;
reg x_reg_L0_22__retimed_I7521_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7521_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296;
	end
assign N13523 = x_reg_L0_22__retimed_I7521_QOUT;
reg x_reg_L0_22__retimed_I7512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7512_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[12];
	end
assign N13500 = x_reg_L0_22__retimed_I7512_QOUT;
reg x_reg_L0_22__retimed_I7500_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7500_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477;
	end
assign N13466 = x_reg_L0_22__retimed_I7500_QOUT;
reg x_reg_L0_22__retimed_I7499_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7499_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228;
	end
assign N13462 = x_reg_L0_22__retimed_I7499_QOUT;
reg x_reg_L0_22__retimed_I7498_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7498_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950;
	end
assign N13460 = x_reg_L0_22__retimed_I7498_QOUT;
reg x_reg_L0_22__retimed_I7497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7497_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853;
	end
assign N13458 = x_reg_L0_22__retimed_I7497_QOUT;
reg x_reg_L0_22__retimed_I7494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7494_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148;
	end
assign N13448 = x_reg_L0_22__retimed_I7494_QOUT;
reg x_reg_L0_22__retimed_I7489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7489_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139;
	end
assign N13436 = x_reg_L0_22__retimed_I7489_QOUT;
reg x_reg_L0_22__retimed_I7488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7488_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387;
	end
assign N13432 = x_reg_L0_22__retimed_I7488_QOUT;
reg x_reg_L0_22__retimed_I7487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7487_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143;
	end
assign N13430 = x_reg_L0_22__retimed_I7487_QOUT;
reg x_reg_L0_22__retimed_I7485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7485_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215;
	end
assign N13424 = x_reg_L0_22__retimed_I7485_QOUT;
reg x_reg_L0_22__retimed_I7452_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7452_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087;
	end
assign N13337 = x_reg_L0_22__retimed_I7452_QOUT;
reg x_reg_L0_22__retimed_I7451_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7451_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157;
	end
assign N13335 = x_reg_L0_22__retimed_I7451_QOUT;
reg x_reg_L0_22__retimed_I7445_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7445_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361;
	end
assign N13319 = x_reg_L0_22__retimed_I7445_QOUT;
reg x_reg_L0_22__retimed_I7442_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7442_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381;
	end
assign N13311 = x_reg_L0_22__retimed_I7442_QOUT;
reg x_reg_L0_22__retimed_I7440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7440_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305;
	end
assign N13305 = x_reg_L0_22__retimed_I7440_QOUT;
reg x_reg_L1_16__retimed_I7411_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I7411_QOUT <= N11929;
	end
assign N13227 = x_reg_L1_16__retimed_I7411_QOUT;
reg x_reg_L1_16__retimed_I7410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I7410_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854;
	end
assign N13225 = x_reg_L1_16__retimed_I7410_QOUT;
reg x_reg_L0_22__retimed_I7409_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7409_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235;
	end
assign N13222 = x_reg_L0_22__retimed_I7409_QOUT;
reg x_reg_L0_22__retimed_I7408_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7408_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171;
	end
assign N13220 = x_reg_L0_22__retimed_I7408_QOUT;
reg x_reg_L0_22__retimed_I7407_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7407_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303;
	end
assign N13218 = x_reg_L0_22__retimed_I7407_QOUT;
reg x_reg_L0_22__retimed_I7404_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7404_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325;
	end
assign N13209 = x_reg_L0_22__retimed_I7404_QOUT;
reg x_reg_L0_22__retimed_I7403_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7403_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418;
	end
assign N13207 = x_reg_L0_22__retimed_I7403_QOUT;
reg x_reg_L0_22__retimed_I7402_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7402_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948;
	end
assign N13205 = x_reg_L0_22__retimed_I7402_QOUT;
reg x_reg_L0_22__retimed_I7401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7401_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413;
	end
assign N13201 = x_reg_L0_22__retimed_I7401_QOUT;
reg x_reg_L0_22__retimed_I7400_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7400_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514;
	end
assign N13199 = x_reg_L0_22__retimed_I7400_QOUT;
reg x_reg_L0_22__retimed_I7399_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7399_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035;
	end
assign N13197 = x_reg_L0_22__retimed_I7399_QOUT;
reg x_reg_L0_22__retimed_I7396_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7396_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104;
	end
assign N13189 = x_reg_L0_22__retimed_I7396_QOUT;
reg x_reg_L0_22__retimed_I7364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7364_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086;
	end
assign N13104 = x_reg_L0_22__retimed_I7364_QOUT;
reg x_reg_L0_22__retimed_I7360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7360_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478;
	end
assign N13094 = x_reg_L0_22__retimed_I7360_QOUT;
reg x_reg_L0_22__retimed_I7359_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7359_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021;
	end
assign N13091 = x_reg_L0_22__retimed_I7359_QOUT;
reg x_reg_L0_22__retimed_I7358_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7358_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739;
	end
assign N13089 = x_reg_L0_22__retimed_I7358_QOUT;
reg x_reg_L0_22__retimed_I7357_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7357_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509;
	end
assign N13087 = x_reg_L0_22__retimed_I7357_QOUT;
reg x_reg_L0_22__retimed_I7355_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7355_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278;
	end
assign N13081 = x_reg_L0_22__retimed_I7355_QOUT;
reg x_reg_L0_22__retimed_I7352_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7352_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479;
	end
assign N13074 = x_reg_L0_22__retimed_I7352_QOUT;
reg x_reg_L0_22__retimed_I7327_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7327_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110;
	end
assign N13004 = x_reg_L0_22__retimed_I7327_QOUT;
reg x_reg_L0_22__retimed_I7326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7326_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209;
	end
assign N13002 = x_reg_L0_22__retimed_I7326_QOUT;
reg x_reg_L0_22__retimed_I7325_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7325_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736;
	end
assign N13000 = x_reg_L0_22__retimed_I7325_QOUT;
reg x_reg_L0_22__retimed_I7311_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7311_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480;
	end
assign N12963 = x_reg_L0_22__retimed_I7311_QOUT;
reg x_reg_L0_22__retimed_I7287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7287_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831;
	end
assign N12897 = x_reg_L0_22__retimed_I7287_QOUT;
reg x_reg_L0_22__retimed_I7286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7286_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297;
	end
assign N12895 = x_reg_L0_22__retimed_I7286_QOUT;
reg x_reg_L0_22__retimed_I7285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7285_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315;
	end
assign N12893 = x_reg_L0_22__retimed_I7285_QOUT;
reg x_reg_L0_22__retimed_I7282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7282_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481;
	end
assign N12885 = x_reg_L0_22__retimed_I7282_QOUT;
reg x_reg_L0_22__retimed_I7261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029;
	end
assign N12827 = x_reg_L0_22__retimed_I7261_QOUT;
reg x_reg_L0_22__retimed_I7260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017;
	end
assign N12825 = x_reg_L0_22__retimed_I7260_QOUT;
reg x_reg_L0_22__retimed_I7259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517;
	end
assign N12823 = x_reg_L0_22__retimed_I7259_QOUT;
reg x_reg_L0_22__retimed_I7253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482;
	end
assign N12807 = x_reg_L0_22__retimed_I7253_QOUT;
reg x_reg_L0_22__retimed_I7234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7234_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101;
	end
assign N12753 = x_reg_L0_22__retimed_I7234_QOUT;
reg x_reg_L0_22__retimed_I7232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7232_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855;
	end
assign N12748 = x_reg_L0_22__retimed_I7232_QOUT;
reg x_reg_L0_22__retimed_I7231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7231_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218;
	end
assign N12746 = x_reg_L0_22__retimed_I7231_QOUT;
reg x_reg_L0_22__retimed_I7230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7230_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343;
	end
assign N12744 = x_reg_L0_22__retimed_I7230_QOUT;
reg x_reg_L0_22__retimed_I7225_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7225_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483;
	end
assign N12731 = x_reg_L0_22__retimed_I7225_QOUT;
reg x_reg_L0_22__retimed_I7205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7205_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167;
	end
assign N12673 = x_reg_L0_22__retimed_I7205_QOUT;
reg x_reg_L0_22__retimed_I7204_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7204_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041;
	end
assign N12671 = x_reg_L0_22__retimed_I7204_QOUT;
reg x_reg_L0_22__retimed_I7203_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7203_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792;
	end
assign N12669 = x_reg_L0_22__retimed_I7203_QOUT;
reg x_reg_L0_22__retimed_I7195_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7195_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484;
	end
assign N12647 = x_reg_L0_22__retimed_I7195_QOUT;
reg x_reg_L0_22__retimed_I7182_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7182_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103;
	end
assign N12609 = x_reg_L0_22__retimed_I7182_QOUT;
reg x_reg_L0_22__retimed_I7181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7181_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358;
	end
assign N12607 = x_reg_L0_22__retimed_I7181_QOUT;
reg x_reg_L0_22__retimed_I7180_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7180_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732;
	end
assign N12605 = x_reg_L0_22__retimed_I7180_QOUT;
reg x_reg_L0_22__retimed_I7178_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7178_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234;
	end
assign N12599 = x_reg_L0_22__retimed_I7178_QOUT;
reg x_reg_L0_22__retimed_I7173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7173_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485;
	end
assign N12586 = x_reg_L0_22__retimed_I7173_QOUT;
reg x_reg_L0_22__retimed_I7156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7156_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486;
	end
assign N12538 = x_reg_L0_22__retimed_I7156_QOUT;
reg x_reg_L0_22__retimed_I7131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7131_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[26];
	end
assign N12466 = x_reg_L0_22__retimed_I7131_QOUT;
reg x_reg_L0_22__retimed_I7130_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7130_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[26];
	end
assign N12464 = x_reg_L0_22__retimed_I7130_QOUT;
reg x_reg_L0_22__retimed_I7129_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7129_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[25];
	end
assign N12460 = x_reg_L0_22__retimed_I7129_QOUT;
reg x_reg_L0_22__retimed_I7125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7125_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487;
	end
assign N12450 = x_reg_L0_22__retimed_I7125_QOUT;
reg x_reg_L0_22__retimed_I7114_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7114_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488;
	end
assign N12418 = x_reg_L0_22__retimed_I7114_QOUT;
reg x_reg_L0_22__retimed_I7104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7104_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416;
	end
assign N12388 = x_reg_L0_22__retimed_I7104_QOUT;
reg x_reg_L0_22__retimed_I7103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7103_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489;
	end
assign N12386 = x_reg_L0_22__retimed_I7103_QOUT;
reg x_reg_L0_22__retimed_I7093_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7093_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946;
	end
assign N12356 = x_reg_L0_22__retimed_I7093_QOUT;
reg x_reg_L0_22__retimed_I7092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7092_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490;
	end
assign N12354 = x_reg_L0_22__retimed_I7092_QOUT;
reg x_reg_L0_22__retimed_I7080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7080_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548;
	end
assign N12320 = x_reg_L0_22__retimed_I7080_QOUT;
reg x_reg_L0_22__retimed_I7073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7073_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570;
	end
assign N12298 = x_reg_L0_22__retimed_I7073_QOUT;
reg x_reg_L0_22__retimed_I7071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7071_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474;
	end
assign N12294 = x_reg_L0_22__retimed_I7071_QOUT;
reg x_reg_L0_22__retimed_I7064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7064_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478;
	end
assign N12272 = x_reg_L0_22__retimed_I7064_QOUT;
reg x_reg_L0_22__retimed_I7063_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7063_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479;
	end
assign N12270 = x_reg_L0_22__retimed_I7063_QOUT;
reg x_reg_L0_22__retimed_I7062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7062_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996;
	end
assign N12268 = x_reg_L0_22__retimed_I7062_QOUT;
reg x_reg_L0_22__retimed_I7040_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7040_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001;
	end
assign N12206 = x_reg_L0_22__retimed_I7040_QOUT;
reg x_reg_L0_22__retimed_I7036_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7036_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532;
	end
assign N12196 = x_reg_L0_22__retimed_I7036_QOUT;
reg x_reg_L0_22__retimed_I7035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7035_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798;
	end
assign N12194 = x_reg_L0_22__retimed_I7035_QOUT;
reg x_reg_L1_22__retimed_I7032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7032_QOUT <= N12156;
	end
assign N12186 = x_reg_L1_22__retimed_I7032_QOUT;
reg x_reg_L1_22__retimed_I7031_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7031_QOUT <= N12154;
	end
assign N12184 = x_reg_L1_22__retimed_I7031_QOUT;
reg x_reg_L0_22__retimed_I7029_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7029_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931;
	end
assign N12178 = x_reg_L0_22__retimed_I7029_QOUT;
reg x_reg_L0_22__retimed_I7028_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7028_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581;
	end
assign N12176 = x_reg_L0_22__retimed_I7028_QOUT;
reg x_reg_L1_22__retimed_I7025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7025_QOUT <= N12138;
	end
assign N12168 = x_reg_L1_22__retimed_I7025_QOUT;
reg x_reg_L1_22__retimed_I7024_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7024_QOUT <= N12136;
	end
assign N12166 = x_reg_L1_22__retimed_I7024_QOUT;
reg x_reg_L0_22__retimed_I7020_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7020_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722;
	end
assign N12156 = x_reg_L0_22__retimed_I7020_QOUT;
reg x_reg_L0_22__retimed_I7019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7019_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982;
	end
assign N12154 = x_reg_L0_22__retimed_I7019_QOUT;
reg x_reg_L1_22__retimed_I7016_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7016_QOUT <= N12120;
	end
assign N12146 = x_reg_L1_22__retimed_I7016_QOUT;
reg x_reg_L1_22__retimed_I7015_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7015_QOUT <= N12118;
	end
assign N12144 = x_reg_L1_22__retimed_I7015_QOUT;
reg x_reg_L0_22__retimed_I7013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7013_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514;
	end
assign N12138 = x_reg_L0_22__retimed_I7013_QOUT;
reg x_reg_L0_22__retimed_I7012_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7012_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775;
	end
assign N12136 = x_reg_L0_22__retimed_I7012_QOUT;
reg x_reg_L0_22__retimed_I7006_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7006_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484;
	end
assign N12120 = x_reg_L0_22__retimed_I7006_QOUT;
reg x_reg_L0_22__retimed_I7005_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7005_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911;
	end
assign N12118 = x_reg_L0_22__retimed_I7005_QOUT;
reg x_reg_L1_22__retimed_I7003_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7003_QOUT <= N12067;
	end
assign N12112 = x_reg_L1_22__retimed_I7003_QOUT;
reg x_reg_L1_22__retimed_I7002_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7002_QOUT <= N12065;
	end
assign N12110 = x_reg_L1_22__retimed_I7002_QOUT;
reg x_reg_L1_17__retimed_I6997_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I6997_QOUT <= N11924;
	end
assign N12097 = x_reg_L1_17__retimed_I6997_QOUT;
reg x_reg_L1_17__retimed_I6996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I6996_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692;
	end
assign N12095 = x_reg_L1_17__retimed_I6996_QOUT;
reg x_reg_L1_18__retimed_I6995_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I6995_QOUT <= N11919;
	end
assign N12092 = x_reg_L1_18__retimed_I6995_QOUT;
reg x_reg_L1_19__retimed_I6993_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I6993_QOUT <= N11914;
	end
assign N12087 = x_reg_L1_19__retimed_I6993_QOUT;
reg x_reg_L1_20__retimed_I6991_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I6991_QOUT <= N11909;
	end
assign N12082 = x_reg_L1_20__retimed_I6991_QOUT;
reg x_reg_L1_21__retimed_I6989_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6989_QOUT <= N11904;
	end
assign N12077 = x_reg_L1_21__retimed_I6989_QOUT;
reg x_reg_L1_22__retimed_I6987_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6987_QOUT <= N11899;
	end
assign N12072 = x_reg_L1_22__retimed_I6987_QOUT;
reg x_reg_L0_22__retimed_I6985_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6985_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755;
	end
assign N12067 = x_reg_L0_22__retimed_I6985_QOUT;
reg x_reg_L0_22__retimed_I6984_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6984_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491;
	end
assign N12065 = x_reg_L0_22__retimed_I6984_QOUT;
reg x_reg_L1_22__retimed_I6962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6962_QOUT <= N11738;
	end
assign N12014 = x_reg_L1_22__retimed_I6962_QOUT;
reg x_reg_L1_22__retimed_I6961_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I6961_QOUT <= N11736;
	end
assign N12012 = x_reg_L1_22__retimed_I6961_QOUT;
reg x_reg_L0_16__retimed_I6928_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I6928_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993;
	end
assign N11929 = x_reg_L0_16__retimed_I6928_QOUT;
reg x_reg_L0_17__retimed_I6926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I6926_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654;
	end
assign N11924 = x_reg_L0_17__retimed_I6926_QOUT;
reg x_reg_L0_18__retimed_I6924_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I6924_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924;
	end
assign N11919 = x_reg_L0_18__retimed_I6924_QOUT;
reg x_reg_L0_19__retimed_I6922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I6922_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572;
	end
assign N11914 = x_reg_L0_19__retimed_I6922_QOUT;
reg x_reg_L0_20__retimed_I6920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I6920_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962;
	end
assign N11909 = x_reg_L0_20__retimed_I6920_QOUT;
reg x_reg_L0_21__retimed_I6918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6918_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505;
	end
assign N11904 = x_reg_L0_21__retimed_I6918_QOUT;
reg x_reg_L0_22__retimed_I6916_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6916_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765;
	end
assign N11899 = x_reg_L0_22__retimed_I6916_QOUT;
reg x_reg_L0_22__retimed_I6847_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6847_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29;
	end
assign N11738 = x_reg_L0_22__retimed_I6847_QOUT;
reg x_reg_L0_22__retimed_I6846_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6846_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67;
	end
assign N11736 = x_reg_L0_22__retimed_I6846_QOUT;
INVX3 float_div_cynw_cm_float_rcp_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353), .A(a_exp[7]), .B(a_exp[0]));
AND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I2 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL float_div_cynw_cm_float_rcp_E8_M23_4_I3 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575), .A(a_exp[6]), .B(a_exp[5]), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2355));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I4 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2353), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11575));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I5 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I6 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I8 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I9 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2376), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2395), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2384), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2404));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I10 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I11 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2389));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I12 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .A(a_man[18]), .B(a_man[17]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I13 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I14 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402), .AN(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B(a_man[16]), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2408), .D(a_man[15]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I15 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2393), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2402));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I16 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2387), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2378));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I17 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29), .AN(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I18 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I19 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A(a_man[21]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_4_I20 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A(a_man[20]));
CLKINVX4 float_div_cynw_cm_float_rcp_E8_M23_4_I21 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A(a_man[19]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_4_I22 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I23 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .A(a_man[17]), .B(a_man[16]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I24 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .A(a_man[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I25 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .A(a_man[16]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I26 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I27 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I28 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I29 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I30 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I31 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I32 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3456), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4009), .B1(a_man[20]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I33 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .A(a_man[16]), .B(a_man[17]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I34 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I35 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I36 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I37 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3847), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3627), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I38 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3807), .B1(a_man[21]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I39 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I40 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I41 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I42 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I43 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4020), .B0(a_man[19]), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I44 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052), .A(a_man[19]), .B(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I45 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I46 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I47 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I48 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3250), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4010), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I49 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3821), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3413), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I50 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I51 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I52 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013), .A(a_man[17]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I53 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I54 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3666), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3280), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I55 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I56 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I57 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3827), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I58 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3414), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4005), .B1(a_man[21]));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I59 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .A1N(a_man[19]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I60 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I61 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I62 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3455), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3281), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I63 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4021), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3624), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I64 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I65 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7962), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7825), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7987));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I66 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I67 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I68 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3502));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I69 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3625), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I70 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I71 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I72 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3356), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I73 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I74 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3294), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3824), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I75 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N499));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I76 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I77 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7505), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7491), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7755));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I78 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I79 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I80 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I81 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I82 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I83 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I84 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3251), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I85 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I86 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I87 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3273), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I88 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I89 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I90 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I91 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3647), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3416), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I92 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3944), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3605), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I93 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I94 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I95 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3820), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3361), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I96 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I97 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I98 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I99 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3848), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3979), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3812), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3620), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3211), .B1(a_man[22]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .A0(a_man[16]), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3980), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3609), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3438), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3214), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3743), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3396), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3618), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4092), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3651), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3648), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3779), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3610), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3408), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3943), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I131 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686), .A(1'B1), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N498));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7572), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7911), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7484));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7639));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .A(a_man[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3375), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3398), .B1(a_man[20]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3233), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3946), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3539), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4131), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3406), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3885), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3443), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3439), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3574), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3399), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3208), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3742), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I166 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17]), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3587), .A1N(a_man[21]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .A(a_man[14]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .A(a_man[13]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4052));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741), .B(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3527), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4117), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16]), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3604));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I178 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6059), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6085));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I179 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[33]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6466), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6524));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I180 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N495), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[33]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I181 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7556));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I182 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7848), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7696), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7686));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4108), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4133), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3601), .B0(a_man[18]), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3966), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3335), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3930), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3205), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3686), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3236), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3234), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3374), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4134), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3942), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3538), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .A(a_man[12]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3561), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3321), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3913), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3846), .B(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3394), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3526), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I215 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6520), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6577));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .A(a_man[11]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3359), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3917), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3748), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4047), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3708), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3926), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4090), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4120), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4130), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3320), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I231 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6114), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6198));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I234 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6480), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6547), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6068));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I235 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[32]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6335), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6255), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5771));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I236 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[32]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[32]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I237 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N494), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7634));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I238 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7453), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7770), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7785));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7654), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7982), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7722));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4123), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3927), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3900), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3933), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3765), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3862), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4061), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3727), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3937), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3478), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3968), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3558), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4107), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3934), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3740), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3334), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .A(a_man[10]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3713), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I272 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3843), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3506), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I273 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3985), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3741), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3883), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3918), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3928), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4046), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I280 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6574), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5823));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I281 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6171), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6141), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6324));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[14]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I286 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5766), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5738), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5796));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I287 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5838), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6289), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5805));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I288 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[31]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6446), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5993), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6369));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I289 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[31]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[31]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I290 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N493), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7716));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I291 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7798), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7665), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7843), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7887));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3329), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3698), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3729), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3557), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3663), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3860), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3523), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3293), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3738), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3271), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3767), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4087), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3899), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3730), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3537), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4060), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .A(a_man[9]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I318 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I319 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3884), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3510), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3340), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3644), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3298), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I324 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I325 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I326 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I327 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3521), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3786), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I328 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3870), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3982), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3684), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3714), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3725), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3842), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I333 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6168), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6308));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I337 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6223), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6196), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6250));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I338 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6135), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5790), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6163));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .A(a_man[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I342 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5763), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5793));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[13]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I345 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5742), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6279), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6463));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I346 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6544), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6512), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6026));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I347 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[30]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6180), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6212), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5729));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I348 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[30]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[30]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I349 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7478), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N492), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7791));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I350 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7532), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8001), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7878), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7927), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7980));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I351 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736), .A(N12194), .B(N12196));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3514), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3495), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3529), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3357), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3453), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3661), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3318), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3535), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4000), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I371 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3564), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3881), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3697), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3530), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3332), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3859), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .A(a_man[7]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I384 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3477), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4029), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I390 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3866), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3559), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I391 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3230), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3826), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I392 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I393 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4038), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3379), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3460), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3577), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3268), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3304), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3316), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3434), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I404 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6221), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6419));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[12]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I407 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6185), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5905));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3685), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3303), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4068), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3766), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3435), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4025), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I421 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3314), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3580), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I422 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .B0(a_man[18]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3671), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3781), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3476), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3511), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3522), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3643), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I428 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5821), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5932), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5848));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I429 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6494), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6117), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5978));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I433 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6248), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6306));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .A(a_man[6]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I439 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3269), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3832), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3393), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3667), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3358), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3963), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3626), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I446 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I447 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3428), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4113), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3256), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3378), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3998), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4031), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4041), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3229), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I456 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5818), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6039));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I458 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6336), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6245), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6364));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I459 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6559), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6416), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6072));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I460 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6008), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6356), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5867));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I461 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[29]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6403), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6054), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6432));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I462 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7996), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[29]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[29]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I463 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7479), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7570), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N491), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7873));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I464 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605), .A(N12270), .B(N12268), .CI(N12272));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3286), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3322), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I471 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I472 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3235), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I475 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I476 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4086), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3247), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3452), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4043), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I481 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B(a_man[18]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3253), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3328), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3803), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I486 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3703), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3363), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3682), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I490 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3323), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N490), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4059), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3660), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I495 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I497 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5873), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5846), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5902));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I498 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5997), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6395), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5760));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I499 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6305), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5930), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6451));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[10]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I502 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I503 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .A(a_man[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I504 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I505 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I506 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4053), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I507 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3999), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3631), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3753), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3457), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4088), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3762), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3415), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3825));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3954), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3906), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3242), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3986), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4111), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3801), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3833), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3839), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3962), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I525 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6274), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6532));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I526 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I527 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6015), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5935), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5931));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I530 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5987), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5959), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6056));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I531 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6373), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6138), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6515));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I532 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5820), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5963), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6195));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I533 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[28]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6243), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6388), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5897));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I534 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7474), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7946), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[28]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[28]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I535 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676), .A(N12354), .B(N12356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I536 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7690), .B(N12294), .CI(N12298));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3655), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I541 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I543 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4016), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4048), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3880), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3977), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3245), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3840), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I548 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I552 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4076), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4055), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3597), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4093), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3474), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3285), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4049), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N489), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3857), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3451), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I566 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6417), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6502), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6447));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I567 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5949), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6201), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6327));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I571 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6333), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6302), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6361));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .A(a_man[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I573 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .A(a_man[3]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I578 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I579 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3596), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3217), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I580 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I581 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I582 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3981), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3683), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3353), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3945), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I588 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3547), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3500), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I592 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4039), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3670), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3582), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3702), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3389), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3423), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3553), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I601 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6331), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5778));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I605 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5906), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6069), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6125));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I606 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I608 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3909), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3395), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I612 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3802), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3421), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I613 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I614 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3905), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4074), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3252), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3882), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3554), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3213), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3828), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3754), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3704), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3788), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3904), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3595), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3632), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3638), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3761), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I630 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5871), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6151));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I632 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6475), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6107), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6392));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I633 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6121), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6001), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6498));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I637 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5928), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5898), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5956));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I640 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I641 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5985), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6095), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6012));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I642 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6487), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5744), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6378));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I643 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5825), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6310), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6434));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I644 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5732), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6087), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6579), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5840));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I645 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6407), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5775), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5917));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I646 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6259), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5883), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6028));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I647 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[27]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5852), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6340), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6573));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I648 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7548), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7416), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[27]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[27]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I649 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776), .A(N12386), .B(N12388));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I650 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7903), .B(N12320), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7676));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I654 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3817), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3844), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3360), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3681), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3776), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3640), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3853), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3390), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I666 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3533), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3688), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3265), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3845), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N488), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3659), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3244), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I671 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I675 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6390), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6359), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6414));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I676 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5921), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6037), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6281));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I677 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I679 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I680 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6443), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6556), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6473));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .A(a_man[2]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .A(a_man[0]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .A(a_man[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I687 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6387));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I688 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5927), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6096));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I690 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6529), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6192), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5726));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I691 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6172), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5798), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6295));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I692 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6011), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5888), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6264));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I693 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I696 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6499), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5747), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5723));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I697 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6188), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6549), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5812));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I698 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5792), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5780), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6391), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5901));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6103), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6216), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6469), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5981));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I700 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[26]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6292), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6148), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6528));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I701 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500), .A(N12464), .B(N12466));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I702 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881), .A(N12418), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7500));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I703 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7503), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7624), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7776));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3324));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I706 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3400), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I707 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3465));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I708 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I710 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I711 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I713 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2800), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2820), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2600));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I719 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I720 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2681), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2842), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2704));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I721 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2852), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2830), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2706));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I723 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I725 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I726 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2771), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2886), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2711));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I728 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2747), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2783), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2638));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I729 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I730 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I733 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2745), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2722), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2694));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I736 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I737 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I738 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I739 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2803), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2815), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2878));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2642), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2630), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2869));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I741 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2674), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2649), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2791));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I742 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I746 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2670), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2790), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2767));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I750 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I751 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2659), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2734), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2828));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I752 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2632), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2893), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2773));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I753 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2686), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2581), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2717));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I757 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I758 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2593), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2597), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2624));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I759 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2883), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2713), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2699));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I760 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2591), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2801), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2617));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I765 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2775), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2701), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2811));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I766 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I770 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I773 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2784), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2666), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2635));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I774 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2781), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2679), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2735));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I775 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2644), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2797), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2614));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I781 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2779), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2712), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2602));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I782 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2752), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2844), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2655));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I783 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2671), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2853), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2843));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I786 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I787 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2824), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2838));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2884), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2789));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I790 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2719), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2611), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2708));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I791 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2724), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2587), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2879));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I792 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2753), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2786), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2604));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I795 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I796 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I798 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2709), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2691));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I799 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2819), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2850), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2805));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I800 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I801 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I802 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I803 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2647), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2741), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2643));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I804 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2677), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2858), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2665));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I805 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2695), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2864), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2683));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I808 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I810 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2833), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2673), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2829));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I811 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2619), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2650), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2793));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I812 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2826), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2809), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2623));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I813 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I814 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I815 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I816 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2787), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2877));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I817 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I818 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I819 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I820 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2685), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2891), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2680));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I821 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2730), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2885), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2702));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I822 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2759), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2608), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2749));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I826 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2715), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2732));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I827 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I828 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2788), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2855), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2818));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I829 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2845), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2871), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2688));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I833 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I834 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I835 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2609), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2595));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I836 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2867), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2861), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2684));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I837 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2633), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2605), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2774));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I839 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I842 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2727), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2578), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2721));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I843 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2832), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2714), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2854));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I844 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I847 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2585), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2778));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I848 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2615), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2726), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2754));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I850 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I851 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I852 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2616), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2636));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I854 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2769), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2590), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2656));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I855 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I856 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I857 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I860 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2629), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2821));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I861 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2770), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2762), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2626));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I862 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I863 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I864 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I865 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I866 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2807), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2675));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I868 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I869 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_4_I870 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2763), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2894), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2814), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2738));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I872 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2813), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2881));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I873 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2586), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2628), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2839));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I874 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2723), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2868), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2697), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2841));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I875 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2799));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2862), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2744), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2796));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2682), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2621), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2865), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2577));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I878 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2645), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2672));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2731), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2846), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2661));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I880 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2742), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2592));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I881 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2874), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2798), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2806));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I882 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2836));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2689), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2576), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2620));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2583), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2890));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2837), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2817), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I886 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2766));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I887 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2584));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2840), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2831));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I889 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2720));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I890 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2895), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2740));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I891 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2860));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I892 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2816), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2658));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I893 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2678));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I894 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2729), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2757));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I895 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2827));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I896 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2834), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2857));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I897 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2641));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2823), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2606));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I899 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2782));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I900 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2888), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2777));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I901 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2599));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I902 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2596), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2848));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2737));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2733), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2663));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I905 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2880));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2808));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I907 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2802), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2696));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_4_I908 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2588), .AN(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2847), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174), .A(N13822), .B(N13824));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[24]), .A(N12599), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3672), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3341), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I913 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I914 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3404), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3436), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3223), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I918 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I919 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I920 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3264), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3372), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I921 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3226), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I923 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3726), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I924 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I925 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3447), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3924), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I927 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I928 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I929 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I930 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3272), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3798), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I931 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3614), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3437), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I932 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N486), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3243), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3774), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I933 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I934 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3864), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3571), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I935 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I936 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3796), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I937 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I938 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3259), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3590), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I939 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N457));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152), .A(N14513), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5101), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2810), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2768));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217), .A(N12599), .B(N12753));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I943 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339), .A(N14513), .B(N12753));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2634), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2625));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070), .A(N12599), .B(N14505));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I947 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I948 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3751), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3709), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3308), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I950 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3916), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3371), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I951 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915), .A(a_man[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I952 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3989), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3915), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I953 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N456));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I954 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272), .A(N13104), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I955 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5339), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5070), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5272));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I956 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5152), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5217), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5347));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I957 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[24]), .B(N12538), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[24]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I959 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3615), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3645), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I963 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I964 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I965 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I966 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3473), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3572), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I967 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3775), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3432), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I968 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3929), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3579), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3654), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4127), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3872), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3546), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I974 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3479), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3995), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I975 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3816), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3646), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N487), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3449), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3975), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I979 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I980 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6122), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6010), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6181));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3993));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I983 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I984 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I985 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4126), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3949), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3780), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3475), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4083), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3744), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3427), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I992 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I993 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3487), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3290), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I997 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3498), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4125), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3218), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3224), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3352), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1001 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1003 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5954), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6262), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5983));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1004 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1005 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1006 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1007 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6036), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6149), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6065));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1008 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6080), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6566), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6459));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1009 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1010 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1011 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1012 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1013 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6233), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6207), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6091));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1014 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5971), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6093), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6472));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1015 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6563), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6061), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6437));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1018 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6495), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5745), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6526));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1020 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1021 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1023 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5833), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5806), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6553));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1024 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6382), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5877), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6251));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1026 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330), .A(a_man[16]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1030 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3291), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3718), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3543), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1033 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3483), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1034 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1035 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3377), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3996), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1036 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3678), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3336), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3392), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3636), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3313), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3871), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3407), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1040 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3808), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3955), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1043 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1045 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3907), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4018), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1046 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3717), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3747), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1047 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3756), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3876), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1050 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1051 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6376), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5980), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5920));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1054 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6491), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5724), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1055 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5892), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6365), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6267));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1056 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5872), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5861), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6234));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1057 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1058 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1059 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1060 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1061 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4023), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3997), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1062 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3923), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3746), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1063 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4096), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1067 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3576), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3266), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1068 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3877), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3540), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1069 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3520));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1072 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4075), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3619), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1073 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4006), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1077 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1078 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4114), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3289), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1079 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3922), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3950), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1080 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3957), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4082), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1081 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1082 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6412), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5886), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5912));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1086 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6032), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6007), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6063));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1087 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1088 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1089 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1090 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1091 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6178), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6319), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1092 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6284), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6385), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5894));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1096 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1097 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6090), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6346), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6119));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1098 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1099 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1101 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6260), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6204), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6288));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1105 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6471), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6440), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5858));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1106 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6270), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5788), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5801));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1107 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5767), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5784), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6143));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1108 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6003), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6477), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5988));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6348), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5984), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6362));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1110 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6517), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5749), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6247), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5764));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6041), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5855), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5967), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6329), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5842));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1112 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6343), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5952), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6076), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6454));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1113 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6358), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6167), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6275), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6153), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6534));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1114 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[23]), .A(N12671), .B(N12669), .CI(N12673));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1115 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[25]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[24]), .A(N12607), .B(N12605), .CI(N12609));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1116 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[24]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[24]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1117 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7523), .B(N12450), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7783));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1118 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[25]), .B(N12460));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1119 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7713), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7709), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7881));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4097), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3594), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3338), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3275), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3939), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4110), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3799), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3470), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4062), .B1(a_man[21]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3549), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3673), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3206), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3606), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3755), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3889), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3787), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3705), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3819), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3516), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3544), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3550), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3677), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6033));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1144 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6000), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6436), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6467));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1145 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6146), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6405), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6301));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1146 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6161), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6552), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6064));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1147 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6521), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6158), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6537));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1152 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5802), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5970), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5856));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1156 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6523), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6492), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5914));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1160 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6551), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5773), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5829));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1161 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5807), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5915), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6290));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1165 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5884), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5942), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5743));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6182), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6194), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6570));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1167 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6543), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6177), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6051));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1168 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6315), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6031), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6046), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6425));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1169 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6218), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6029), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6139), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6128), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6503));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1170 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[22]), .A(N12746), .B(N12744), .CI(N12748));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1171 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[23]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1172 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7647), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7988), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7859));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1173 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7922), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7568), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7972));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4054), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3804), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3267), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3204), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3231), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3270), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3994), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4104), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3370), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3959), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3947), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3988), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3239), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3719), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3464), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4002), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3592), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3403), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3232), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N485), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3973), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3569), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193), .A(N14513), .B(N14505));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2601), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2812));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258), .A(N12599), .B(N14500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125), .A(N13104), .B(N12753));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1198 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5193), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5258), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5125));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316), .A(N13104), .B(N14505));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385), .A(N14513), .B(N14500));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2703), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2667));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113), .A(N12599), .B(N14510));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1203 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5316), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5385), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5113));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3545), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3575), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3664), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3248), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3450), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3736), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4033), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3711), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4103), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4069));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3508), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N455));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399), .A(N14533), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1215 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5330), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5399), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5169));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5270), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5242), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5390));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1217 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[23]), .B(N12586), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[23]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3343), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3376), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4089), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3534), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3835), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3509), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3895), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3295), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3735), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3536));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3868), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3902), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3586), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3301), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N454));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183), .A(N13081), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247), .A(N14533), .B(N12753));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5171), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2627), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2851));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5303), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5235), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1237 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194), .A(N13220), .B(N13218), .CI(N13222));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1238 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5183), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5247), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5266));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377), .A(N13081), .B(N12753));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5104), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4070), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4109), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3486));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3207), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3327), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3633), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3302), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3694), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4022), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3852), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4013), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3331), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3653), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3668), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3700), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3383), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4027), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N453));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308), .A(N14528), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1257 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5377), .B(N13189), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5308));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1258 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5252), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5077), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5064));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1259 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5315), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5141), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5286));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1260 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1261 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7461), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7730), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7940));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1262 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7526), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7590), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7468));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3274), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3310), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4066), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4004), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1272 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1273 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3903), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3593), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3263), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3861), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3734), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3462), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3940), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3691), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3484), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3581), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3501), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3617), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3309), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3339), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3347), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3469), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1290 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6486), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6060), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6086));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1291 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6213), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5722), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6307));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1292 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6082), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6461), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6557));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1293 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6428), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6442), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5955));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3411), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3983), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4124), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3865), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3603), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3330), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3701), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3387), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3662), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3806), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3637), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3257), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3739), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4132), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3380), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3292), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3405), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4035), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4067), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0]), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4079), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3262), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5990));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1318 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1319 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1321 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5854), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5828), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5998));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1322 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5841), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6175), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6485));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1323 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5994), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6100), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6465));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1324 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5960), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6352), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5864));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1325 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1326 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1327 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1328 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5966), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6578), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5881));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1333 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5741), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6050), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5913));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1334 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5734), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6105), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6118));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1340 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6170), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6199));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1341 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6079), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5769), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6124));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1345 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5939), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6025), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5800));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6401));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1348 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1349 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6374), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6116), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6285));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1350 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6375), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5999), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6496));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1351 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6370), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5979), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6357));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1355 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6144), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6457), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6316));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1359 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6257), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6227), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6404));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1360 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6197), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6575), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5822));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1364 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6344), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6427), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6203));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1365 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5730), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6084), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6481));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1366 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5976), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6070), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6448));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1367 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6509), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6337), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6240), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5753));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1368 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6297), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6110), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6220), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6320), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5834));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1369 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5736), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5944), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6332), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5845));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1370 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6017), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5831), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5938), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6410), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5925));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1371 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[20]), .A(N12895), .B(N12893), .CI(N12897));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3350), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3858), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3733), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3763), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3442), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4030), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3591), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3695), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3893), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3551), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4042), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3584), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1384 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3770), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3311), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3345), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3867), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3461), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3362), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1390 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3600), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4122), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1391 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3935), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3764), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1392 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N483), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3567), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4101), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1393 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[21]), .A(N12825), .B(N12823), .CI(N12827));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1394 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[21]), .B(N12731), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3599), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4077), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3936), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3964), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3446), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3797), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3896), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3758), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3791), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3499), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3970), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3518), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3805), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3386), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3203), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3965), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N484), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3773), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3369), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1414 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[22]), .B(N12647), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1415 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7804), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7753), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7540));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1416 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7734), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7673), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7566));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1418 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6009), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6389), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5899));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1419 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5868), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5880), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6256));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1421 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1422 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1424 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6565), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6225), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6254));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1428 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6513), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6423), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6342));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1429 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5903), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6500), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6294));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1433 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6314), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6283), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6371));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6106), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6548));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1438 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6455), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6484), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6399));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1439 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6516), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6394));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1440 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6261), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5885), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6273));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1441 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6035), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6244), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5772), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6145));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1442 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6209), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6021), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6131), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5849), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6224));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1443 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[19]), .A(N13002), .B(N13000), .CI(N13004));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3307), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4106), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4072), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3417), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1446 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3532), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3555), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1447 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4073), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[18]), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3385), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3491), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3348), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3480), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4019), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3565), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4037), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3792), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3687), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3391), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3920), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3732), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3556), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N482), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3368), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3892), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1463 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[20]), .B(N12807), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[20]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2580), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2892));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2690), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2710));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1469 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5381), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5305), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5345), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5279), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5212));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3524), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1471 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3430), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1472 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3901), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1475 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3941), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1476 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3424), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4028), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3490), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3568), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3793), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3277), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3822), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3566), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1481 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3612), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4057), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3445), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3458), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3497), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4116), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3830), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1486 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092), .A(N14523), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353), .A(N14528), .B(N14505));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079), .A(N13081), .B(N14500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5148), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1490 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5353), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5079), .CI(N13448));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1491 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281), .A(N13311), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5092), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5187));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5087), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5157), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295), .A(N14533), .B(N14500));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1495 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324), .A(N13337), .B(N13335), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5295));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1497 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1498 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1499 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3669), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3699), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3388), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4118), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1502 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3652), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3219), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1503 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3831), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3282), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1504 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1505 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3809), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3790), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1506 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3621), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3365), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1507 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3874), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4056), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3856), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3238), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3254), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3288), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3912), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3629), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N451));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218), .A(N14518), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284), .A(N14523), .B(N12753));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1517 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5215), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5143), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5066), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5337));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1518 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5218), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5284), .CI(N13424));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5361), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229), .A(N13081), .B(N14505));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162), .A(N14528), .B(N12753));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1522 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135), .A(N13319), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5229), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5162));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1523 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5335), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5135));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1524 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5356), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5341), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5165));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1525 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5206), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5398), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5194));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1526 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5374), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5226), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5211));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1527 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[21]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1528 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7612), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7823), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7886));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1529 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7943), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7408), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7668));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1530 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6408), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5918), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1531 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5777), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5791), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6165));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1534 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6022), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6160));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1536 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5922), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6541), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5936));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1540 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6047), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6077), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1541 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1543 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1544 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5910), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5879), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5964));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5945));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1548 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5797), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6104), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5937));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1549 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6190), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5814), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6296));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1550 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6186), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6278), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5795));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1552 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1554 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6136), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5824), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5851));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1555 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5827), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6564), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6202));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1556 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6169), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6561), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6073));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1557 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5948), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6545), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6150), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6530));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1558 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5739), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6413), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6525), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5758), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6137));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1559 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[18]), .A(N13089), .B(N13087), .CI(N13091));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4078), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3326), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3354), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3258), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3634), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3769), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4121), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3283), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3489), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4080), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3750), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3974), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3759), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3440), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1571 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3364), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3837), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3706), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1573 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3585), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3541), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3967), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4128), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3716), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3531), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3355), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N481), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4098), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3692), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1578 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[19]), .B(N12885), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1579 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268), .A(N13081), .B(N14510));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1580 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5139), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1581 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071), .A(N14518), .B(N12753));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1582 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5268), .B(N13436), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5071));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2603), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2751));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5198), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5133), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204), .A(N14528), .B(N14500));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1587 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289), .A(N13601), .B(N13599), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5204));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1588 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5173), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5362), .CI(N13305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5396), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5260), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1592 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3783), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4040), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3459), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3496), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4024), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3548), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3444), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3951), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3630), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4011), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3412), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3492), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3410), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4095), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3349), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3656), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3969), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3984), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4017), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3707), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3419), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1606 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N450));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195), .A(N13725), .B(N12753));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1608 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267), .A(N13557), .B(N13555), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5195));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5122), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2765), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2610));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5389), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1612 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328), .A(N14523), .B(N14500));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1613 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121), .A(N13593), .B(N13591), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5328));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1614 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5343), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5196), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5289));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2748), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2794));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1619 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5223), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5150), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5312), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5240), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5175));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3722), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3990), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3317), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3255), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3287), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3855), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3891), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3382), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4115), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3237), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3749), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3420), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3813), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3528), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3504), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3210), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3209), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3887), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3987));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3921), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3241), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3768), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3784), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3818), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3216), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N449));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127), .A(N13712), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1640 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5370), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5296), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5108), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5382), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5245));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1641 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078), .A(N13549), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5127), .CI(N13551));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340), .A(N13725), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1646 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5387), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5311), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5254), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5189), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5323));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1647 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244), .A(N13430), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5340), .CI(N13432));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1648 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5097), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5155), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5244));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1649 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5073), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5126), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5273));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1650 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5116), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5319), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5261));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1651 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5281), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5147), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5293));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1652 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5102), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5088), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5237));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1653 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5310), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5153), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5297));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1654 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[19]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1655 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7909), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7561));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1656 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[20]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1657 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7543), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7489), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7769));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1661 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6482), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5757));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1665 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6367), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6562), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6398));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1666 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5735), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6094), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6474));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1667 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5721), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6313), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6078));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1671 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6453), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6538), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6309));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1675 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6510), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6339), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6422));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1676 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6363), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5986), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6488));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1677 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6456), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6089), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6470));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1678 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5853), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6452), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6546), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6058));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1679 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6514), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6325), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6038), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6055), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6433));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1680 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[17]), .A(N13199), .B(N13197), .CI(N13201));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3422), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3782), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3402), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4051), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4084), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3623), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3315), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3616), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3919), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4012), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3279), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3873), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1690 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3225), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3658), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1691 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3910), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3737), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1692 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4094), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3635), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1693 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4135), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3854), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3342), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3583), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3560), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1696 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3925), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3513), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1697 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3325), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4085), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1698 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N480), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3890), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3488), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[18]), .B(N12963), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[18]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1700 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7773), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7979), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7427));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1701 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7758), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7959), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7871));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6354));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2887), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1706 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6074), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1707 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5733), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6280), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5787));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1708 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6002), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6109), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5874));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1709 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6246), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5982), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5968), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6360));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1710 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6418), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6228), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6341), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5965), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6435));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1711 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[16]), .A(N13207), .B(N13205), .CI(N13209));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3563), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3578), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1713 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3246), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3851), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3878), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3931), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3715), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3814), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4008), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3675), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1719 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3588), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3777), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3886), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3426), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3503), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3240), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1723 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4001), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3720), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3306), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1725 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4050), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3879), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1726 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N479), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3690), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3278), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1727 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[17]), .B(N13074), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386), .A(N13725), .B(N14505));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1729 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114), .A(N14518), .B(N14500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1730 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5179), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1731 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5386), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5114), .CI(N13709));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318), .A(N13712), .B(N12753));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1733 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2870), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2652));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5234), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1736 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5395), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5320), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5094), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5231));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1737 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1738 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5203), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5130), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5099), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5366), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5299));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1741 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5318), .B(N13689), .CI(N13693));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1742 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228), .A(N13541), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5177), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5304), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5172), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5365));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5164), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1746 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1747 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5378), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5220), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5358));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1748 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084), .A(N13787), .B(N13785), .CI(N13789));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5372), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1750 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5166), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1751 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5236), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1752 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276), .A(N13808), .B(N13806), .CI(N13810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1753 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5161), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5352), .CI(N13659));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1754 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5267), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5121), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5137));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1755 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5393), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5301), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5111));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1756 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5081), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5221), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5368));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1757 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[18]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1758 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7846), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7450), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7512));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1759 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7963), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7637), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7967));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1760 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3562), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4063), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3897), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3650), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3679), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3721), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1765 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3789), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3836), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1766 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3938), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3467), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3512), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3611), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3466), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1770 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3972), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3296), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3689), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3222), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3515), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3220), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3971), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3908), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3800), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3519), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4032), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3850), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3680), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N478), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3485), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4007), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1782 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6101), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5933), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6020));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1783 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1786 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5962), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6156), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5992));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1787 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6540), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5909), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6159));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1790 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1791 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6045), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6132), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6189));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1792 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5799), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6049), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6282));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1793 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6249), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6380), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5765));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1795 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2822), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1796 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6536), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5813));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5895));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1798 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5847), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5904), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6460));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1799 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1800 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1801 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1802 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6420), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5754), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6450));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1803 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1804 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6303));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1806 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6560), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6396), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6479));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1808 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1810 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6507), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5731), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5785));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1811 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6222), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5737), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6113));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1812 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6426), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6174), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5941));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1813 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6535), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6265), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5889), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6140));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1814 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5950), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5762), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5870), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6345), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5857));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[15]), .A(N13460), .B(N13458), .CI(N13462));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1816 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876), .A(N13094), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1817 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1818 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1819 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5342), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5145));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1821 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5144), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5069), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5167), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5089), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5302));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1822 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384), .A(N13675), .B(N13673), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5276));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1823 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5118), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5248), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5400));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5086), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1826 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1827 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5184), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5112), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5224), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5154), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5083));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5158), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5291), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5363), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5292));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1831 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257), .A(N13800), .B(N13798), .CI(N13802));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1832 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232), .A(N13699), .B(N13697), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5332));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1833 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5105), .B(N13523), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5307));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1834 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5283), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5078), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5228));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1835 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[15]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5376), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5090), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5182));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1836 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[16]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1837 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7929), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7876), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7795));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1838 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[16]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5255), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5201), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5349));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1839 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[17]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1840 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7564), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7720), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7459));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741), .A(N13094), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1842 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1843 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1844 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3297), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3731), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3441), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3471), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3367), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3221), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3757), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3911), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3305), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3401), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3607), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3260), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1850 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3333), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4071), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1851 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3823), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4100), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1852 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3481), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3953), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3639), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4034), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3622), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3771), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1855 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3712), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3598), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1856 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3409), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3312), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3834), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1857 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3649), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3472), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N477), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3425), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3276), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3810), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1859 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5974), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6350), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5862));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1860 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6330), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6062), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6550), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6318));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1861 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6231), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6044), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6519), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5782), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6154));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1862 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[14]), .A(N13585), .B(N13583), .CI(N13587));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1863 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477), .A(N13466), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1864 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7741), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7602), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1865 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7778), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7579), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7558));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1868 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1869 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1870 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5123), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5388), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5076), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5214));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1872 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1873 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1874 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5313), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5238), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5346), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5274), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5208));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1875 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216), .A(N13720), .B(N13718), .CI(N13722));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1876 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5290), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5084), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5232));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1877 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[14]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5263), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5207), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5357));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1878 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[15]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7477), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1879 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7984), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7663), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7662));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1880 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1881 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1882 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6130), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6268));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5850));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1886 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6016), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6214), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6040));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1887 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6522), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6287), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5804));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1889 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1890 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1891 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6155), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6187), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6071));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1892 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6411), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6179), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6034));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1893 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6237), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6490), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6005));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1894 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6030), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5844), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5832), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6439), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5953));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1895 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[13]), .A(N13609), .B(N13607), .CI(N13611));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1896 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1897 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1899 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2648), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1900 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5728), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5865));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1901 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6241), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6098), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6242));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1902 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6258));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1905 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5752), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5811), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6501));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1907 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1908 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1909 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6533), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5783), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6558));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1910 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5756), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6099), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6134));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1911 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5926), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6555), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6067));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1912 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6206), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6384), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5751), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6129));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1913 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[12]), .A(N13733), .B(N13731), .CI(N13735));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1914 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5146));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1918 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5249), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5391));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1919 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5062), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5327), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5067), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5199), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5192));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1920 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344), .A(N13771), .B(N13769), .CI(N13773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1921 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1923 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5371), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5129), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5265));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1924 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1925 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5278), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1927 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5178), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5401), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5333));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1928 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5269), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5197), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5091), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5106), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5250));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1929 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5257), .B(N13681), .CI(N13685));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1930 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5216), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5080), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5364));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1931 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[13]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[13]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1932 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5384), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5098), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5190));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1933 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[14]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[14]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1934 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7800), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7861));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1935 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7456));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1936 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7585), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[15]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7762));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1937 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7723));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1938 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1939 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1941 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6184), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2579), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1943 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6572), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5839), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6053));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1944 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6478), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5991), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6511));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1945 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6445), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6300), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5816));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1946 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5893), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6506), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6019));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1947 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1948 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1950 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5338), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5264), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5256), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5185), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5120));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1951 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138), .A(N13880), .B(N13878), .CI(N13882));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1952 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5209), .B(N13630), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5344));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1953 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[12]), .B(N13500), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1954 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8004), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[13]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7961));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1955 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1956 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1959 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6152), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6238), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6293));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5808));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1963 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6211), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6266), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6126));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1964 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6462), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6083), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6431));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1965 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6024), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6368), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5878));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1966 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[10]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5958), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6193), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6569));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1967 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5205), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1968 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1969 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5379), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1971 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5151), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5075), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5085), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5325), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5119));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1972 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[10]), .A(N13763), .B(N13761), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5138));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1973 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550), .A(N13649), .B(N13647), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[11]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1974 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7452), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7607), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[12]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1975 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1979 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5809), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5863), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5836));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1982 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5779), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5919));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1983 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5929), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6415), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6386));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1984 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5977), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5946), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6322));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1985 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[9]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6253), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6402), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5770));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5334));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1989 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5233), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5110), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5309), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5241));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1990 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[9]), .A(N13872), .B(N13870), .CI(N13874));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1991 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651), .A(N13779), .B(N13777), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1992 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7819), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7550));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1993 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6215));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1997 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1998 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6232), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6381));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1999 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5890), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5748), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5774));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2000 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6304), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5896), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6271));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2001 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5837), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6355), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6210));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5132), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2003 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5259));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2004 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5163), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5300));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2005 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2006 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5397), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5186));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2009 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5287), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5156));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5367), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5095), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5321));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5354), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5131), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5277));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2012 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757), .A(N13864), .B(N13862), .CI(N13866));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2013 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7423), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[10]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7651));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2014 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2018 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6263), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6323), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6291));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6226), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6147), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5740));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2020 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[8]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5789), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5819), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6162));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2021 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851), .A(N13898), .B(N13896), .CI(N13900));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2022 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[9]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7757));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2023 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2024 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2026 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5916), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2028 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6372), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6351), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6449));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2029 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[7]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6115), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6527), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6493));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2030 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7839), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7949), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[7]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2031 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974), .A(N13837), .B(N13835), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7851));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2033 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6166));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2034 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2035 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2036 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5859), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5887), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5975));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2037 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[6]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5961), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5882), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6338));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2039 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7445), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2040 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574), .A(N13890), .B(N13888), .CI(N13892));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5115));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2043 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2045 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6377), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6406));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2046 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2875), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2047 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6576));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6120));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2050 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5969), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6027));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2051 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6430), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6347), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6102));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2052 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[5]), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6183), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6483), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5996));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5322), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2054 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2055 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7925), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7789), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7656), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7444));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969), .A(N13842), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2057 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5246), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N5380));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2058 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2059 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7528), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7868), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7546));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2060 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711), .A(N13854), .B(N13856));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2061 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7642));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2062 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2063 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[3]));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2066 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[2]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2067 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2068 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6568), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6531), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6299), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N6075));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2069 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7895), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7414));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7547), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7811));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7525), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7636), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7990));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2072 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7786), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7487), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7945), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7597));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2073 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7737), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7995));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7623), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7436), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7857), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7921));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7711), .A1(N13852), .B0(N13854), .B1(N13856));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831), .A(N13842), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7574));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2077 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7969), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7926), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7831));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2078 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7625), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7609), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7715), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7974));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2079 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7506), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7767));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2080 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7902), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7828), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7763));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2081 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7549), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7442), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7905), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7555));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7693), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7951));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7814), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7583), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7688));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7476), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7733), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7481), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7745));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7882), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7534));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7739), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7796), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7599));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2087 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7997), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7860), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7667), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7933));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2088 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22792), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7694), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22794), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N22796));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2089 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2090 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7552), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N11605), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7852), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7515));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7641), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7912), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7431), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7701));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7827), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7492), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2096 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7619), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7891));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2097 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2098 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7412), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7678), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2099 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7808), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7465));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7595), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7865), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7992), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7652));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7440), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7787), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7571), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7835));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7971), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7628), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7764), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7420));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593), .A0N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7551), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7817), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7605), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7948));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467), .A(N12206), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415), .A0N(N12206), .A1N(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7742), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510), .B1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415), .B0(N12194), .B1(N12196));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7993), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7581), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7931));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7692), .A0N(N12176), .A1N(N12178), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7854), .B1(N11929));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438), .A0(N12097), .A1(N12095), .B0(N12184), .B1(N12186));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7924), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7775), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7514));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806), .A0N(N12166), .A1N(N12168), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438), .B1(N12092));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486), .A0(N12087), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806), .B0(N12144), .B1(N12146));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768), .AN(N12082), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486));
OA22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970), .A0(N12077), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768), .B0(N12110), .B1(N12112));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7614));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N4112), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3952));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N3894), .B(a_man[22]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7765), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7889), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7790));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[39]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7970), .B(N12072));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I2132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2523), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2514), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2526), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2518));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2516), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7]), .A(a_exp[7]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5]), .A(a_exp[5]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3]), .A(a_exp[3]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1]), .A(a_exp[1]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[0]), .A(a_exp[0]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2139 (.CO(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464), .S(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2]), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2459));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2457));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2451));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_4_I2149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3]), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6]), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2449));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4]), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2464));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483), .AN(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2489), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4]), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2486), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2483));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17), .A0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[7]), .A1(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N2444), .B0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N446));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__9));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33), .AN(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N447), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34), .D(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I2161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__67), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N448));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2162 (.Y(x[22]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[39]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[38]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7768), .B(N12077));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2164 (.Y(x[21]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[38]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[37]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7486), .B(N12082));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2166 (.Y(x[20]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[37]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[36]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7806), .B(N12087));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2168 (.Y(x[19]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[36]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[35]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7438), .B(N12092));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2170 (.Y(x[18]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[35]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[34]), .A(N12095), .B(N12097));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2172 (.Y(x[17]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[34]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[33]), .A(N13225), .B(N13227));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2174 (.Y(x[16]), .A(N12014), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[33]), .S0(N12012));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7415), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7736));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[15]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[32]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7510), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7467));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[14]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[31]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7593), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7809));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[13]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[30]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7604), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7544));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[12]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[29]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7618), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7893));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[11]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[28]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7554), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7620));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[10]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[27]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7495), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7964));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[9]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[26]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7954), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7703));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[8]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[25]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7812), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7432));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[7]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[24]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7592), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7779));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[6]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[23]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7978), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7517));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[5]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[22]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7689), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7853));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[4]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[21]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7991), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7586));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[3]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[20]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7617), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7934));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[2]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[19]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7850), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N7669));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[1]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[18]), .S0(N11736));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8002), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_N8005));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[0]), .A(N11738), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[17]), .S0(N11736));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_4_I2208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__34), .C(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__33));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[7]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[6]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[5]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[4]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[3]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[2]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2215 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[1]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2216 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__42));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[31]), .AN(a_sign), .B(float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__29));
reg x_reg_L0_23__I2241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__I2241_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[23];
	end
assign N5603 = x_reg_L0_23__I2241_QOUT;
reg x_reg_L0_24__I2242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_24__I2242_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[24];
	end
assign N5608 = x_reg_L0_24__I2242_QOUT;
reg x_reg_L0_25__I2243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_25__I2243_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[25];
	end
assign N5613 = x_reg_L0_25__I2243_QOUT;
reg x_reg_L0_26__I2244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_26__I2244_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[26];
	end
assign N5618 = x_reg_L0_26__I2244_QOUT;
reg x_reg_L0_27__I2245_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_27__I2245_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[27];
	end
assign N5623 = x_reg_L0_27__I2245_QOUT;
reg x_reg_L0_28__I2246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_28__I2246_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[28];
	end
assign N5628 = x_reg_L0_28__I2246_QOUT;
reg x_reg_L0_29__I2247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__I2247_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[29];
	end
assign N5633 = x_reg_L0_29__I2247_QOUT;
reg x_reg_L0_30__I2248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_30__I2248_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[30];
	end
assign N5638 = x_reg_L0_30__I2248_QOUT;
reg x_reg_L0_31__I2249_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I2249_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[31];
	end
assign N5643 = x_reg_L0_31__I2249_QOUT;
reg x_reg_L1_0__I2250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__I2250_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[0];
	end
assign x[0] = x_reg_L1_0__I2250_QOUT;
reg x_reg_L1_1__I2251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__I2251_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[1];
	end
assign x[1] = x_reg_L1_1__I2251_QOUT;
reg x_reg_L1_2__I2252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__I2252_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[2];
	end
assign x[2] = x_reg_L1_2__I2252_QOUT;
reg x_reg_L1_3__I2253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__I2253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[3];
	end
assign x[3] = x_reg_L1_3__I2253_QOUT;
reg x_reg_L1_4__I2254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__I2254_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[4];
	end
assign x[4] = x_reg_L1_4__I2254_QOUT;
reg x_reg_L1_5__I2255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__I2255_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[5];
	end
assign x[5] = x_reg_L1_5__I2255_QOUT;
reg x_reg_L1_6__I2256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__I2256_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[6];
	end
assign x[6] = x_reg_L1_6__I2256_QOUT;
reg x_reg_L1_7__I2257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__I2257_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[7];
	end
assign x[7] = x_reg_L1_7__I2257_QOUT;
reg x_reg_L1_8__I2258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__I2258_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[8];
	end
assign x[8] = x_reg_L1_8__I2258_QOUT;
reg x_reg_L1_9__I2259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__I2259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[9];
	end
assign x[9] = x_reg_L1_9__I2259_QOUT;
reg x_reg_L1_10__I2260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__I2260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[10];
	end
assign x[10] = x_reg_L1_10__I2260_QOUT;
reg x_reg_L1_11__I2261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__I2261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[11];
	end
assign x[11] = x_reg_L1_11__I2261_QOUT;
reg x_reg_L1_12__I2262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__I2262_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[12];
	end
assign x[12] = x_reg_L1_12__I2262_QOUT;
reg x_reg_L1_13__I2263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__I2263_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[13];
	end
assign x[13] = x_reg_L1_13__I2263_QOUT;
reg x_reg_L1_14__I2264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__I2264_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[14];
	end
assign x[14] = x_reg_L1_14__I2264_QOUT;
reg x_reg_L1_15__I2265_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__I2265_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[15];
	end
assign x[15] = x_reg_L1_15__I2265_QOUT;
reg x_reg_L1_23__I2273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__I2273_QOUT <= N5603;
	end
assign x[23] = x_reg_L1_23__I2273_QOUT;
reg x_reg_L1_24__I2274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__I2274_QOUT <= N5608;
	end
assign x[24] = x_reg_L1_24__I2274_QOUT;
reg x_reg_L1_25__I2275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__I2275_QOUT <= N5613;
	end
assign x[25] = x_reg_L1_25__I2275_QOUT;
reg x_reg_L1_26__I2276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__I2276_QOUT <= N5618;
	end
assign x[26] = x_reg_L1_26__I2276_QOUT;
reg x_reg_L1_27__I2277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__I2277_QOUT <= N5623;
	end
assign x[27] = x_reg_L1_27__I2277_QOUT;
reg x_reg_L1_28__I2278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__I2278_QOUT <= N5628;
	end
assign x[28] = x_reg_L1_28__I2278_QOUT;
reg x_reg_L1_29__I2279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__I2279_QOUT <= N5633;
	end
assign x[29] = x_reg_L1_29__I2279_QOUT;
reg x_reg_L1_30__I2280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__I2280_QOUT <= N5638;
	end
assign x[30] = x_reg_L1_30__I2280_QOUT;
reg x_reg_L1_31__I2281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I2281_QOUT <= N5643;
	end
assign x[31] = x_reg_L1_31__I2281_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__22[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_2_inst_inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  srLwTgzZqxw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



