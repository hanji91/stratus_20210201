/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:06:45 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_2 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42;
wire [15:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710,
	float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737;
wire N12256,N12258,N12260,N12465,N12467,N12472,N12474 
	,N12479,N12481,N12486,N12488,N12493,N12495,N12500,N12502 
	,N12547,N12549,N12569,N12762,N12772,N12782,N12784,N13010 
	,N13012,N13026,N13085,N13189,N13191,N13310,N13375,N13432 
	,N13440,N13450,N13460,N13470,N13480,N13490,N13500,N13502 
	,N13517,N13519,N13521,N13537,N13539,N13547,N13549,N13551 
	,N13557,N13559,N13561,N13584,N13586,N13588,N13592,N13594 
	,N13596,N13600,N13602,N13604,N13608,N13610,N13612,N13616 
	,N13618,N13620,N13624,N13626,N13628,N13632,N13634,N13636 
	,N13640,N13642,N13644,N13648,N13650,N13652,N13666,N13668 
	,N13670,N13673,N13678,N13680,N13682,N13693,N13695,N13697 
	,N13715,N13717,N14033,N14061,N14065,N14304,N14305,N14306 
	,N14307,N14308,N14309;
reg x_reg_19__retimed_I8143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I8143_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589;
	end
assign N14065 = x_reg_19__retimed_I8143_QOUT;
reg x_reg_14__retimed_I8141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I8141_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746;
	end
assign N14061 = x_reg_14__retimed_I8141_QOUT;
reg x_reg_14__retimed_I8128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I8128_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960;
	end
assign N14033 = x_reg_14__retimed_I8128_QOUT;
reg x_reg_15__retimed_I8010_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I8010_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848;
	end
assign N13717 = x_reg_15__retimed_I8010_QOUT;
reg x_reg_15__retimed_I8009_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I8009_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690;
	end
assign N13715 = x_reg_15__retimed_I8009_QOUT;
reg x_reg_2__retimed_I8000_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I8000_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770;
	end
assign N13697 = x_reg_2__retimed_I8000_QOUT;
reg x_reg_2__retimed_I7999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7999_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[11];
	end
assign N13695 = x_reg_2__retimed_I7999_QOUT;
reg x_reg_2__retimed_I7998_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7998_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[11];
	end
assign N13693 = x_reg_2__retimed_I7998_QOUT;
reg x_reg_2__retimed_I7995_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7995_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579;
	end
assign N13682 = x_reg_2__retimed_I7995_QOUT;
reg x_reg_2__retimed_I7994_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7994_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283;
	end
assign N13680 = x_reg_2__retimed_I7994_QOUT;
reg x_reg_2__retimed_I7993_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7993_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130;
	end
assign N13678 = x_reg_2__retimed_I7993_QOUT;
reg x_reg_2__retimed_I7991_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7991_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607;
	end
assign N13673 = x_reg_2__retimed_I7991_QOUT;
reg x_reg_2__retimed_I7990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7990_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683;
	end
assign N13670 = x_reg_2__retimed_I7990_QOUT;
reg x_reg_2__retimed_I7989_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7989_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[12];
	end
assign N13668 = x_reg_2__retimed_I7989_QOUT;
reg x_reg_2__retimed_I7988_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7988_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946;
	end
assign N13666 = x_reg_2__retimed_I7988_QOUT;
reg x_reg_2__retimed_I7984_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7984_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213;
	end
assign N13652 = x_reg_2__retimed_I7984_QOUT;
reg x_reg_2__retimed_I7983_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7983_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203;
	end
assign N13650 = x_reg_2__retimed_I7983_QOUT;
reg x_reg_2__retimed_I7982_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7982_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222;
	end
assign N13648 = x_reg_2__retimed_I7982_QOUT;
reg x_reg_18__retimed_I7981_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7981_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[18];
	end
assign N13644 = x_reg_18__retimed_I7981_QOUT;
reg x_reg_18__retimed_I7980_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7980_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[18];
	end
assign N13642 = x_reg_18__retimed_I7980_QOUT;
reg x_reg_18__retimed_I7979_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7979_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928;
	end
assign N13640 = x_reg_18__retimed_I7979_QOUT;
reg x_reg_2__retimed_I7978_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7978_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206;
	end
assign N13636 = x_reg_2__retimed_I7978_QOUT;
reg x_reg_2__retimed_I7977_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7977_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214;
	end
assign N13634 = x_reg_2__retimed_I7977_QOUT;
reg x_reg_2__retimed_I7976_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7976_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233;
	end
assign N13632 = x_reg_2__retimed_I7976_QOUT;
reg x_reg_15__retimed_I7975_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7975_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282;
	end
assign N13628 = x_reg_15__retimed_I7975_QOUT;
reg x_reg_15__retimed_I7974_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7974_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[20];
	end
assign N13626 = x_reg_15__retimed_I7974_QOUT;
reg x_reg_15__retimed_I7973_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7973_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[20];
	end
assign N13624 = x_reg_15__retimed_I7973_QOUT;
reg x_reg_15__retimed_I7972_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7972_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098;
	end
assign N13620 = x_reg_15__retimed_I7972_QOUT;
reg x_reg_15__retimed_I7971_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7971_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[21];
	end
assign N13618 = x_reg_15__retimed_I7971_QOUT;
reg x_reg_15__retimed_I7970_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7970_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[21];
	end
assign N13616 = x_reg_15__retimed_I7970_QOUT;
reg x_reg_15__retimed_I7969_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7969_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294;
	end
assign N13612 = x_reg_15__retimed_I7969_QOUT;
reg x_reg_15__retimed_I7968_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7968_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[22];
	end
assign N13610 = x_reg_15__retimed_I7968_QOUT;
reg x_reg_15__retimed_I7967_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7967_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[22];
	end
assign N13608 = x_reg_15__retimed_I7967_QOUT;
reg x_reg_18__retimed_I7966_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7966_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733;
	end
assign N13604 = x_reg_18__retimed_I7966_QOUT;
reg x_reg_18__retimed_I7965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7965_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[19];
	end
assign N13602 = x_reg_18__retimed_I7965_QOUT;
reg x_reg_18__retimed_I7964_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7964_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[19];
	end
assign N13600 = x_reg_18__retimed_I7964_QOUT;
reg x_reg_2__retimed_I7963_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7963_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243;
	end
assign N13596 = x_reg_2__retimed_I7963_QOUT;
reg x_reg_2__retimed_I7962_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7962_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230;
	end
assign N13594 = x_reg_2__retimed_I7962_QOUT;
reg x_reg_2__retimed_I7961_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7961_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225;
	end
assign N13592 = x_reg_2__retimed_I7961_QOUT;
reg x_reg_2__retimed_I7960_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7960_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575;
	end
assign N13588 = x_reg_2__retimed_I7960_QOUT;
reg x_reg_2__retimed_I7959_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7959_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[13];
	end
assign N13586 = x_reg_2__retimed_I7959_QOUT;
reg x_reg_2__retimed_I7958_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7958_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835;
	end
assign N13584 = x_reg_2__retimed_I7958_QOUT;
reg x_reg_15__retimed_I7950_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7950_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862;
	end
assign N13561 = x_reg_15__retimed_I7950_QOUT;
reg x_reg_15__retimed_I7949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7949_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221;
	end
assign N13559 = x_reg_15__retimed_I7949_QOUT;
reg x_reg_15__retimed_I7948_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7948_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[26];
	end
assign N13557 = x_reg_15__retimed_I7948_QOUT;
reg x_reg_15__retimed_I7947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7947_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664;
	end
assign N13551 = x_reg_15__retimed_I7947_QOUT;
reg x_reg_15__retimed_I7946_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7946_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054;
	end
assign N13549 = x_reg_15__retimed_I7946_QOUT;
reg x_reg_15__retimed_I7945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7945_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[25];
	end
assign N13547 = x_reg_15__retimed_I7945_QOUT;
reg x_reg_15__retimed_I7943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7943_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267;
	end
assign N13539 = x_reg_15__retimed_I7943_QOUT;
reg x_reg_15__retimed_I7942_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7942_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244;
	end
assign N13537 = x_reg_15__retimed_I7942_QOUT;
reg x_reg_2__retimed_I7937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7937_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236;
	end
assign N13521 = x_reg_2__retimed_I7937_QOUT;
reg x_reg_2__retimed_I7936_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7936_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[14];
	end
assign N13519 = x_reg_2__retimed_I7936_QOUT;
reg x_reg_2__retimed_I7935_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7935_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747;
	end
assign N13517 = x_reg_2__retimed_I7935_QOUT;
reg x_reg_2__retimed_I7930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7930_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[15];
	end
assign N13502 = x_reg_2__retimed_I7930_QOUT;
reg x_reg_2__retimed_I7929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7929_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657;
	end
assign N13500 = x_reg_2__retimed_I7929_QOUT;
reg x_reg_15__retimed_I7926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7926_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718;
	end
assign N13490 = x_reg_15__retimed_I7926_QOUT;
reg x_reg_15__retimed_I7923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7923_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745;
	end
assign N13480 = x_reg_15__retimed_I7923_QOUT;
reg x_reg_18__retimed_I7920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7920_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128;
	end
assign N13470 = x_reg_18__retimed_I7920_QOUT;
reg x_reg_2__retimed_I7917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7917_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198;
	end
assign N13460 = x_reg_2__retimed_I7917_QOUT;
reg x_reg_15__retimed_I7914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7914_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942;
	end
assign N13450 = x_reg_15__retimed_I7914_QOUT;
reg x_reg_2__retimed_I7911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I7911_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211;
	end
assign N13440 = x_reg_2__retimed_I7911_QOUT;
reg x_reg_15__retimed_I7909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7909_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913;
	end
assign N13432 = x_reg_15__retimed_I7909_QOUT;
reg x_reg_18__retimed_I7890_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7890_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307;
	end
assign N13375 = x_reg_18__retimed_I7890_QOUT;
reg x_reg_11__retimed_I7871_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7871_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003;
	end
assign N13310 = x_reg_11__retimed_I7871_QOUT;
reg x_reg_14__retimed_I7830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7830_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630;
	end
assign N13191 = x_reg_14__retimed_I7830_QOUT;
reg x_reg_14__retimed_I7829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7829_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214;
	end
assign N13189 = x_reg_14__retimed_I7829_QOUT;
reg x_reg_19__retimed_I7796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7796_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185;
	end
assign N13085 = x_reg_19__retimed_I7796_QOUT;
reg x_reg_14__retimed_I7777_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I7777_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783;
	end
assign N13026 = x_reg_14__retimed_I7777_QOUT;
reg x_reg_19__retimed_I7772_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7772_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768;
	end
assign N13012 = x_reg_19__retimed_I7772_QOUT;
reg x_reg_19__retimed_I7771_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7771_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604;
	end
assign N13010 = x_reg_19__retimed_I7771_QOUT;
reg x_reg_11__retimed_I7690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7690_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889;
	end
assign N12784 = x_reg_11__retimed_I7690_QOUT;
reg x_reg_11__retimed_I7689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I7689_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047;
	end
assign N12782 = x_reg_11__retimed_I7689_QOUT;
reg x_reg_12__retimed_I7685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I7685_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008;
	end
assign N12772 = x_reg_12__retimed_I7685_QOUT;
reg x_reg_13__retimed_I7681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I7681_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198;
	end
assign N12762 = x_reg_13__retimed_I7681_QOUT;
reg x_reg_19__retimed_I7607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I7607_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692;
	end
assign N12569 = x_reg_19__retimed_I7607_QOUT;
reg x_reg_15__retimed_I7599_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7599_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170;
	end
assign N12549 = x_reg_15__retimed_I7599_QOUT;
reg x_reg_15__retimed_I7598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I7598_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737;
	end
assign N12547 = x_reg_15__retimed_I7598_QOUT;
reg x_reg_22__retimed_I7579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7579_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817;
	end
assign N12502 = x_reg_22__retimed_I7579_QOUT;
reg x_reg_22__retimed_I7578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7578_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989;
	end
assign N12500 = x_reg_22__retimed_I7578_QOUT;
reg x_reg_21__retimed_I7576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I7576_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080;
	end
assign N12495 = x_reg_21__retimed_I7576_QOUT;
reg x_reg_21__retimed_I7575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I7575_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242;
	end
assign N12493 = x_reg_21__retimed_I7575_QOUT;
reg x_reg_20__retimed_I7573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I7573_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584;
	end
assign N12488 = x_reg_20__retimed_I7573_QOUT;
reg x_reg_20__retimed_I7572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I7572_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752;
	end
assign N12486 = x_reg_20__retimed_I7572_QOUT;
reg x_reg_18__retimed_I7570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7570_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846;
	end
assign N12481 = x_reg_18__retimed_I7570_QOUT;
reg x_reg_18__retimed_I7569_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7569_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015;
	end
assign N12479 = x_reg_18__retimed_I7569_QOUT;
reg x_reg_17__retimed_I7567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I7567_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108;
	end
assign N12474 = x_reg_17__retimed_I7567_QOUT;
reg x_reg_17__retimed_I7566_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I7566_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265;
	end
assign N12472 = x_reg_17__retimed_I7566_QOUT;
reg x_reg_16__retimed_I7564_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I7564_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616;
	end
assign N12467 = x_reg_16__retimed_I7564_QOUT;
reg x_reg_16__retimed_I7563_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I7563_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774;
	end
assign N12465 = x_reg_16__retimed_I7563_QOUT;
reg x_reg_18__retimed_I7472_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7472_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67;
	end
assign N12260 = x_reg_18__retimed_I7472_QOUT;
assign N14304 = !N12260;
assign N14305 = !N14304;
reg x_reg_18__retimed_I7471_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7471_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934;
	end
assign N12258 = x_reg_18__retimed_I7471_QOUT;
assign N14306 = !N12258;
assign N14307 = !N14306;
reg x_reg_18__retimed_I7470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I7470_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320;
	end
assign N12256 = x_reg_18__retimed_I7470_QOUT;
assign N14308 = !N12256;
assign N14309 = !N14308;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127 = !(a_exp[6] & a_exp[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813 = !((a_exp[7] & a_exp[0]) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3125);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3127 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13813);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 = !a_man[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167 = !((((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142) | a_man[0]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3163) | a_man[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161 = !(((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3148 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3169) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3158) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3179);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0] = !((((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3167) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3161) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3173) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3183);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328 = !(((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3326) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3338) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3330);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3328 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1] = !a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0] = !a_exp[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2] = !a_exp[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2] = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3] = !a_exp[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3240) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5] = !a_exp[5];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4] = !a_exp[4];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[3] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3256 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3246);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5] = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5] ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3248;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[5] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6] = !a_exp[6];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3241));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3254 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7] = !a_exp[7];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3233) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3244);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0] = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[0] ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[4];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3250) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289 = !((((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3295) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[8] = !((((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3247) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[6]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3237) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__20[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3289 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3292) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[8];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3209 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__17);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__30) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__9 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3320 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N447;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688 = ((float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[0]) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26688;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9934 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__67;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 = !a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 = !a_man[21];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 = !a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350 = !a_man[18];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 = !a_man[20];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4350;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 = !a_man[16];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4601 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5015;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516 = !a_man[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13759;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4385 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4246 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4821 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4867 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4979 | a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N501;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141 = !(a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4646 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4231 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4468 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4824 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4374 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5025 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 = !(a_man[17] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4418 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4232 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5042 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4600 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N500;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4419 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5029 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4847 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4603 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4156 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4803 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5041 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[19] & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4198 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5030 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4817 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4373 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N499;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4516 & a_man[16]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 & a_man[17]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4421;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4199 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4225 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4626 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4376 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4955 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4581 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4816 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4319 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4848 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4993 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4808 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4596 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4155 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976} = {1'B0, 1'B1} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N497};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9133 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8771);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8948 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8749 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9147);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9129 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9240)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8989 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8909;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8817 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9234 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8957;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4206) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 = !(a_man[17] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13767;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4713;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4994 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4585 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13789;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4400 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4158 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4728 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4358 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & a_man[17]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4594 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5117 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4631 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4627 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4770 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4586 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4369 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4954 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] = !a_man[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4334 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4360 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13748;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4180 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4957 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4508 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5157 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13558;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4367 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4890 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13761;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4613 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4825;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4405 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4401 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4546 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4361 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4152 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4727 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N495};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N496) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9192;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4495 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5143 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16] = !(a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4580);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 = !a_man[14];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4560 & a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 = !a_man[13];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7205} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[17]);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[33], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[32]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7595} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7656} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4777 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5133 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5160 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4576 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4980 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4292 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4938 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4149 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4669 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4183 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4181 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4333 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5161 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4952 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4507 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[32]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[33]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9026} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8631};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 = !a_man[12];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4532 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4275 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4920 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4926 | a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4356 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4494 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15]);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7651} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7710};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4934 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5115 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5145 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4317 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4924 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4734 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5069 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4691 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4274 & a_man[22]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5156));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 = !a_man[11];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7233} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7322} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[16];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7680} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7609} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7188};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[32], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[31]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7380} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7463} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6882};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5148 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4935 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4906 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4941 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4862 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5083 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4709 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4947 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4445 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4982 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4529 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5132 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4942 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4724 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4291 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[31]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9218} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[32]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8814};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 = !a_man[10];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7707} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6849} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7261} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7293} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7451};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4705 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5001));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4726 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4888) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4925 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826) ^ a_man[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5116 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4695));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4844 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4473 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645 = !((a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5068) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4936));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7339;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6935} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6877} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6908};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7415} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6950} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6917};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[31], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[30]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7112} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7573} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7498};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4285 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4681 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4711 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4528 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4643 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4860 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4492 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4245 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4722 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4223 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4756 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5112 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4905 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4712 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4506 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5082 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[30]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8662} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[31]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9014};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8768 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 = !a_man[9];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7290} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4889 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4477));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4298) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4622 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (a_man[21] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4251));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4490 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4778 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4873) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4997 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4667 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (a_man[21] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4696));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[12] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4707 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4843 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[12];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7435} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7347} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7375};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6902} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7254} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7285};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 = !a_man[8];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6874} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6905} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7645;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7405} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6853} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7591};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7642} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7676} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7147};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[30], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[29]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7336} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7301} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6840};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4482 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4461 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4497 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4315 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4416 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4641 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4272 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4504 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5019 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4536 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4886 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4680 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4498 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4288 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4859 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[29]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[30]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9207};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4444) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5051));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4868 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4530 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4176 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4823 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5059 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4338));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4424 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4549 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4220 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4257 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4269 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4396 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7547} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7402} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7432};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7067;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4668) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4256));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5091 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4755 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4397 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5047 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4267 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4552 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4651 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4772 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4443 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4478 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4491 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4621 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7464} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7523};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7544} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7693} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7192};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 = !a_man[7];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7373} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6990} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7022} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7307};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[11]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7051} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6933} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6961};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 = !a_man[6];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6929} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6958} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4221 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4830));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5081 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4647 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4316 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4975 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4602 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4391 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5138 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4205 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4337 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5017 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5053 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5063 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4175 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7160} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6988} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7019};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7370} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6871};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7048} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7431} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7579};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7128} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7516};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7236} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7624} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7097};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[29], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[28]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7560} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7530};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4238 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4277 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4182 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5111 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4196 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4415 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5066 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4202 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4284 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4798 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4687 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4321 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4664 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4460 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4278 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5080 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4640 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[10];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7049} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7136} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7078};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 = !a_man[5];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7399} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7054} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7176};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7258} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7646};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6932} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7318};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[28], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[27]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6981} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7013} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7368};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[28]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[29]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9039} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8648};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8589 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4636 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13762 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5036 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5070 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4885 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4991 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4193 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4841 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5100 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5077 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4571 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5118 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4441 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4237 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5071 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4858 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4414 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[27]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[28]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9231} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8830};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4591 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4623 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4440 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4544 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4765 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4394 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4937 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4635 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5152 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4877 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4446 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5013 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4812 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4624 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4412 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4989 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4299 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4365 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4398 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4215 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4330 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4542 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4173 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13764 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4708 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4551 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4410 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4932 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4224 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4792 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4590 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4399 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4191 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4764 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5076 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4799 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4148 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4178 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4995 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4222 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5012 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5129 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4328 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4972 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4958 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5005 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4187 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4702 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5021 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4565 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4364 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4179 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4987 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4541 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4573 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4945 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4977 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4902 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5126 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4746 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4784 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4465 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4984 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4486 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4800 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4347 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4147 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4978 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4763 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4327 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4308 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4716 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4752 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4404 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5052 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4564 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4678 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4899 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4522 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4264 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13763 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4303 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4425 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4320 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4574 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5147 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4944 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4753 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4539 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5125 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4260 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5131 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5096 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4500 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4526 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5097) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4346 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4456 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4676 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4306 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5007;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5040 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4537 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5058 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4353 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4928 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4715 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4527 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4326 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4898 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4282 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4312 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4818 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4759 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5146 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4235 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4454 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5104 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4988 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4322 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4836 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4558 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4510 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5153 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4698 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4499 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4313 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5123 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4675 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4382 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4773 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4363 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5073 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5109 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4927 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5032 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4230 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4878 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4172 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4917 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5119 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4612 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4855 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4556 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4933 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4481 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4281 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5110 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4895 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4453 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4534 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4629 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4661 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4835 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4480 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4588 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4807 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4430 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4986 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4249 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4672 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4168 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4985 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4915) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4487 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5054 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4850 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4662 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4451 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5027 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4535 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4851 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4883 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4411 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4697 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4810 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5028 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4657 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4971 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13807 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4891 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4388 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4188 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5020 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4703 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4259 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5072 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4884 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4673 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4229 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N479};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8588};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N481} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9157};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8970};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8767};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8574};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N485} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9142};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8953};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N487} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8754};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4409 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4813 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4845 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4318 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4663 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4767 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4990 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4618 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4854 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4352 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4900));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4501 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4671 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4216 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5035 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4846 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4639 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4192 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4916) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4740));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4357) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4797 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4381 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4912 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5098 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4201 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4887 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4525 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4157 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4742 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4688));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4431));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4780 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4910));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4569 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (a_man[21] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4608));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4617) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4749));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4670 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5075 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5022));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5018 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4607 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4741) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4420 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5113 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4750 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4375 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4822);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4966) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4913));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4190 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5002 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5137));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4796 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4831 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4839 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4974 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7271} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7046} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7244};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7075} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7105} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7133};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6856} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7616} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7121};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7068} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7712};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 = !a_man[4];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6986} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7014} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 = !a_man[3];
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7458} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7487} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4177 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4170 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4570 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4163));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4969 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4428 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4652 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4592 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4996 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4665 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4311 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4956 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4517 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13791 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4518 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4466));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5060 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4650 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4554 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4686 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4351 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4383 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4393 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4524));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6891} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7518} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6837};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7023} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7039} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7407};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7545} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7574} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7227};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7571} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7661} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7602};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[7];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[9];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7542} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6859} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7690};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6910} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7294} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7422};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7005} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7388};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7157};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5010);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5064));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5151 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4961 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4771) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4442 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5107) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4729 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4470 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4390));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4452 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4304 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4242));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4903 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4340 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4464 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5150 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4164 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4171 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4310));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5]);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7045} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7386};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7630} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6834};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6923} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7311} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7682};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[8]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7664} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7460} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7489};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7520} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7633} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7604};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7507} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7629};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7519} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6893} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7018};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7598} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7340} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7101};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7437} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6937} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7325};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7000} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7149} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7383};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7454} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7208} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6953};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7535} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7035};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[26], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[25]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7268} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7419} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7660};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8862} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8893} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[26]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[27], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[26]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7468} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6964} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7706};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9003} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[27]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9029} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8675};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9047 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695 = !(N13191 & N12782);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156 = !(N14065 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030 = !(N13012 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4279);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4439 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 = a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4429;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571 | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3683} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3661} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3421};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3499 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3669);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3723) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3676} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3750} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3664};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3414} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3418} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3716};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3648} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3501} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3620};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13732} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3487} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3690};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3758} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3558} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3542};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3774} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3454} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3626};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3663} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3444};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3569} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3596} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3537};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3453} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3467} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3743};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3397} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3564};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3544} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3672} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3422};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3498} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3458} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3646};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26325} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26352};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3656} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3470} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3437};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3556} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3634} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3630};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3450} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3601} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3482};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3725} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3715};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3765} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3625} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3554};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3474} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3510} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3649};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3713} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3518} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3548};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3637} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3461};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3692} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3550};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3687} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3706};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3571;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3591} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3473};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26335} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26340} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26307};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26322} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26349} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26318};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3640} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3604} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3425};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3759) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3638;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3553} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3535};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3682} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3468} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3666};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26338} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26333};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26341};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3641} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3749};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3772} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3729} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3525};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3761} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3547};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3691} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3698} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3507};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26327} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26314};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3612} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3433} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3598};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26363} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26359} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26330};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3434} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3416};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26598};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3562} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3583};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3517} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3681};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3428} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3628};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3744} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3718} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3532};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3395} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3577};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26621} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26601} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26626};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3402} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3633};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26583} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26603} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26608};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3441} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3460};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26610} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26593};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26629 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26634);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | (!a_man[7]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3452} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3685};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3615} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3623} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3451};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26637;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26615;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | (!a_man[6]));
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3668} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3511};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3617) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3555)) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3674) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3588));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3624 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3404) | (!(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3673 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3754)));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3570) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3526)) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3541) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3712));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26616 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26624);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26638) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26619 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26611);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26606 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26627) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26587 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26579));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26590 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26596;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26581) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26636)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3593 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3413);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3753 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3621) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3540);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3489 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3703);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3400 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3771);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3574 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3710) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3483);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3464 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3619);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3709 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3694);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3775 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3590);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3678 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3486);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3580 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3609);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3700 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3731);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3429 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3686);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3767 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3632);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3417 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3719);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3584 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3494);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424 = !(((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3708)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3618));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3500)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3424);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3699) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3608);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3549)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3459);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3546) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3629);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[24] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3488 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3411));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3705) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3466;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4964);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4864 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4543 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4563 & a_man[22]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4209);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3717 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3627));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3403);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3480 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3704 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3737);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3600 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3582;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3463);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3565 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3530;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3475) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3512)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3430);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3768) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3419)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3720);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3528) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3442);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3675) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3766)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3684);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3762) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3680);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4738 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4692 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4261 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4923 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4329 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922 = !(a_man[21] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5006 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4922 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N456;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6385} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6182} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6451};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[24], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6264} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6329} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6459};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8586} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[24]};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7130} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7331} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7269};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 = !a_man[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 = !a_man[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7515};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7073} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7217} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7103};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7302} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7156} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7241};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7700} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7200} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7587};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[6];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7359} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7212};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7091} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7214} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7601};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7181} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7697} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7566};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6918} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6857};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[5];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4981 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5045 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5016 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4931) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4732));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4869 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5121 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4785 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4548) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4217 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4882 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (a_man[21] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4509));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4489);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5099 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4595 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5026) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4218 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5139 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4241 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4930 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4962 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[4] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4970 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5106 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[4];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7540} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6971} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7003};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7606} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7108} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7123};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7600} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6888} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6835};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6945} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7028} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7658};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6992} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7510};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7104} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6974};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7071} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7582};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7274} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7401} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7666};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[25], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[24]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7223};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9221, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9054} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8731} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[25]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193} = {1'B0, N13557} + {1'B0, N13559} + {1'B0, N13561};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600 & N13310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4550 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4243 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4701 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4512 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4449 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4336 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5014 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4660 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4293 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4354) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4615));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4266));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4876 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4368));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4804) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4967));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4914 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5039 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4700 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4733 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[3] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4744 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4881));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7505} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7038};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7625} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7686} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7621};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7009} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7391};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7360} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6987};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7183} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7153} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7356};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7127} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7384};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7414} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7328} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7238};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7513} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7011} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7394};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6896} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6878} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7279};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7372} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6861} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6875};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7456} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7087} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6955};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[24], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6904} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7162} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7289};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8664, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9244} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8925} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[24]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634} = {1'B0, N13547} + {1'B0, N13549} + {1'B0, N13551};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5093);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4768));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4515 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4547 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4644 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4968 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4413 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4720 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5055 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4694 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5128 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399 = !((a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26412) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26419));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26399;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3545 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3455));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3670;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3647 | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3751));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3734 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3594;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3506) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3427);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6511} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6305} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6371};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4739 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5101 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4706 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4301 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4335 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4271 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4503 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4834 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4476 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4901 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4247 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4718 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4505);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4871 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4908 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4559 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4254 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N454;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3760 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3679));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3478) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3560) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3644);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6225} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6295} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6428};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6237} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6442} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6281};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[23], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[22]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6355} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6383} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6502};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9267, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[23]};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6855;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7475} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7299};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6913} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6900} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7410};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7576);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5122 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4402 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4568 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4485 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4295));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4438 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4227) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4949));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4794 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4747));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5136 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4793 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4434 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (a_man[21] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5085));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4721 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4520 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4599));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4654 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4150));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13797) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4582) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4743 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4894 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4689 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4815 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4484 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4513 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4521 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4659));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2]);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7596} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7565} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7120};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7622} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7001} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7031};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7266} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7532} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7032};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7685} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7298} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7283};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7263} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7669} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7652};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7159;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6941} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7090} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6884};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7655} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6969} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6914};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7684} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7061} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6833};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7416} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6919} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7303};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7317} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7428} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7703};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7184} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7675} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7171};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7166} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7152} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7553};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7247} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7634};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[23], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[22]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7472} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7342} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6968};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8848, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8690} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9110} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[23]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818} = {1'B0, N13537} + {1'B0, N13539} + {1'B0, N13717};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4226 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4263 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5089 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5024 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13782 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4166));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4557 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4909 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4566 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4213 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4861 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4194 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4717 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5127 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4427 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4950 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13744);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13760 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4450 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4553 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4467 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4593 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4262 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4296 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4433 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6998);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7180} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7615} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7442};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7503} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7555} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7411};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7433} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6854} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6934};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7202} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7589} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7691};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7570} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7556} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7074};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7206} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7473};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7264} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7235} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7296};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7320} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7708};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7531} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7352};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7204} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7610};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7095} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7575};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7459} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7063} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6957};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7538} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7057} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7043};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[22], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[21]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7648} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7138} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7150};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8718, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9294} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[22]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8980} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[22]};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3592 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3504));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26111;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4584 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4619 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5043 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4852 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5141 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4287 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4633 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4648 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4683 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4377 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5094 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5134 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4151 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5061 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13766 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4610 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4255 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4677 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26095 & a_man[22]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26089 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26100;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6415} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6420};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6360} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6379};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6283} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6489};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6176};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[22], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[21]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6253} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6427} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6399};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881} = {1'B0, N13608} + {1'B0, N13610} + {1'B0, N13612};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017} = {1'B0, N13490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9042} + {1'B0, N13715};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4371 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4998 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5149 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5057 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4865 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4297);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4579 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4286 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4685 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4348 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5009 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4642 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4802 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5102 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4252 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4616 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4208) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4723));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5158 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4561 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4736 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4339));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4244 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (a_man[20] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4366));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5056 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5090 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5103) | (a_man[22] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4212));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[15] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7304);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7681} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7058} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7170};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7327} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6954} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7225};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7221} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7113} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7593};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7481} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6977};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6852} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7029} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6880};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7086} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7711} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6997};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6966} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7117} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6940};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6845} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7614} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7118};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7237} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7129} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7517};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7098} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7499} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7485};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7551} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7349};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6912} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7243};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7626} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7015} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7504};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6982} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6996} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7381};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7465} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6962};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7446} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6946};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[21], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[20]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7441} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7424} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6943};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8913, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8745} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9172} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[21]};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3742 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3662);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[17] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3491) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3426 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3726));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3642;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3747) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3559;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3394) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3509) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3696);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6392} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6324};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13795 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4939 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4435 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4207 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4649 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4682 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5088 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4632 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4165 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4829 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4234 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4875 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13803 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4300 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13772));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4805 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4597 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4323 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4879 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & a_man[17]) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5078 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4857 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4186 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4203 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4240 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4919 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4605 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N451;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6330} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6465};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6274} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6299};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3471 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3392));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3631;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3589 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3579) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3485);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3523) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3439);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6245} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6310};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5108 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4349 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4392 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4872 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4907 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4280 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4953 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13786));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4951 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4783 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4386 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5050 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4455 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4540 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4786) | (a_man[19] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4276));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4819 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4538 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4344 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5079 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4408 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4422 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4463 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5142 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4828 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N452;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6327} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6191} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6397};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6269} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6473} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6199};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6342} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6204} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6407};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6436} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6447} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6247};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6453} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6468} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6277};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6510} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6318} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6306};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[21], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[20]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6339} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6323};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7533);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7292} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7323};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7226) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7146;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7470} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7527} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7583};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7647} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7631} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7522};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3538 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7409} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7699} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7673};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7613} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7500} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7440};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7135} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7020} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7036};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7002} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7398} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7385};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7536} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7421} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6921};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6889} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6903} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7287};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6883} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7369} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6870};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6865} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7348};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[20], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7333} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6847} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7229};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9098, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8942} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8605} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[20]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070} = {1'B0, N13616} + {1'B0, N13618} + {1'B0, N13620};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9235} + {1'B0, N13432} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8881};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5087 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4774 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5062 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4423 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4462 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5046 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4519 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4268 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4948 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4407 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4963 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4606 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5031 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4372 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5124 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4457 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4370 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5120 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4307 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13752 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4637 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4983 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5000 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5037 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4690 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4379 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N450;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6452} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6316};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6449} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6178} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6381};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6474} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6417};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6435} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6367} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6301};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6183} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6255} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6499};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6228} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6431} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6374};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6394} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6405};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[20], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6422} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6409};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7143} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6936};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7040} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7055};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7083} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7056} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6995};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7224} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7197} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7026};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6952);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7114} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7167} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6909};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7423} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6925} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7313};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7404} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7308} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6907};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7270} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7677} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7175};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7657} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7256};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[19], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7639} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6850} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7142};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9282, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9128} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8792} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[19]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257} = {1'B0, N13624} + {1'B0, N13626} + {1'B0, N13628};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653} = {1'B0, N13480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8680} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9070};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4704 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4531 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4162 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4270 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4204 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4239 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4856 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4897 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4341 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5140 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4185 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4735 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4380 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4809 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4496 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4471 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4154 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4153 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4892 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5004);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5163 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4929 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4189 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4758 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4776 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4814 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4472 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4161 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N449;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6286);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6239} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6373} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6440};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3695 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3605));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3730 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3763;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6508} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6501} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6234};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6308} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6455} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6401};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3521 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3438));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3508;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227 = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3659) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3575);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6424} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6353} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6220};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3534 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26096);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26097 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26104);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26090) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26108);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6358} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6287};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6336} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6307} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6482};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6209} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6267} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6357};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6238} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6386};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[19], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6200} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6214} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6350};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3496 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7282} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7255} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6963};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7698} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7439} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7326};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7291} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7695} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7193};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7257);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7611} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7406};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7550} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7526} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7467};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7215} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6846} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7106};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6939} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6832} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7198};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3462 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7640} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6869};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7696} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7670} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7495};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7603} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7228};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7194} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7052};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7436} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6844} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6899};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7617} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7122} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6989};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7210} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7584} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7088};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7679} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7580} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7178};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7662} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7561} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7158};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[18], float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7155} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7644} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7541};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8733, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9307} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8994} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[18]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707} = {1'B0, N13600} + {1'B0, N13602} + {1'B0, N13604};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833} = {1'B0, N13450} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8866} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9257};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6213);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6291} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6498} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6430};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6423} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6233};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6278};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3739 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3657));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6347 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6478} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6206} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6211};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6507} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6226} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6315};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6416} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6411} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6484};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6403} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6470};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6477);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6490} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6349} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6284};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6464} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6262} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6273};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6380} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6438} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6249};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6505} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6413} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6223};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[18], float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26243} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6333} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26266} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6480};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7277} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7081};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7111} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7222};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7025} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7672};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7508} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7006};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7599} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7102} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7474};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7564} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7084} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7469};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26233} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7066} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7546} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7452};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8928, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26198} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26236} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26263};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898} = {1'B0, N13640} + {1'B0, N13642} + {1'B0, N13644};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032} = {1'B0, N13470} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9056} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8707};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3432 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7165} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7312};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7169} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7408} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6911};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6983);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7668} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7524};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7562);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7021} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6960} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7588};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7295} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7554} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7683};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6876} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7389} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7260};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6970} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6985};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26203} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6965} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7069} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7353};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N478;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4314) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13754 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13788));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4656 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4250 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4714 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4403 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4436 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4325 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4167 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4918 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4258 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4362 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4583 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4210 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4290 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5095 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4820 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N5159 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4447 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4965 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13745 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13806) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4479 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4598 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4849 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4533) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4572 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4265 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4896) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4833 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4628 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4634) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4437 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4228 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4911) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N4806 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7608} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7694} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7578};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6866} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6842} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7548};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3399 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7637} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6924} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6897};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7346} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6848} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7232};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7093} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6975};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7060} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7182} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7444};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6894} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7650} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7275};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[15], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7357} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7371} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6873};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26222} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26230, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26214} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8840} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26240};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6276 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6266} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6332} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6337};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6201} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6195} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6270};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6296} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6432} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6444};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6408} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6217} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6419};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6396} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6341};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26225, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26211} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26219} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26246} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26253};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227} = {1'B0, N13592} + {1'B0, N13594} + {1'B0, N13596};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9246} + {1'B0, N13375} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8898};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6404);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6257} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6188};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6279} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6475} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6414};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6242} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6256} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6389};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6361} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6230} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6512};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26206, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[15]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6202} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26229};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247} = {1'B0, N13632} + {1'B0, N13634} + {1'B0, N13636};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667} = {1'B0, N13460} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26227};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6331);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6320} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6393} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6326};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6198 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6387} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6454} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6458};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6425} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6235} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6224};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6402} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6345};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26213, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6469};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7276};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7288);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7338} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7309} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7137};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7413} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7654} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6916};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7191} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7161} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7219};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7300} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7539};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7620} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7362} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7125};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7567} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6944} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7072};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[14], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7151} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7667} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7164};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3702 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6839} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6864};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7392} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7366} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7367};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6922} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6895} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7692};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7594);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3611 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7665} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7632} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6978};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6868} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7253};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7689} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7044} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7187};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6863} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7512} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7248};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[13], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7330} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6956};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6437} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6503};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6304};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6351} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6500};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6378} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6311};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3714);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3756 | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26407));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6467 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26415) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26417);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6513} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6241} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6246};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6218} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6203} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6363};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6370} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6181};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[13], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6192} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6328} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6476};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8747, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8575} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[13]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[14], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6210} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6496} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6302};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8657, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9236} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[14]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807} = {1'B0, N13517} + {1'B0, N13519} + {1'B0, N13521};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720} = {1'B0, N13648} + {1'B0, N13650} + {1'B0, N13652};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562} = {1'B0, N13500} + {1'B0, N13502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8720};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7306} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7335};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7705} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6951} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7173};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7607} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7110} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7641};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7427} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7572} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6927};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[12], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7010} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7636} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7140};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6391 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6184);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6297} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6362} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6369};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6290};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[12], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6321} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6309} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6456};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8835, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8683} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[12]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918} = {1'B0, N13584} + {1'B0, N13586} + {1'B0, N13588};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3446 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7016);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7245} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7453} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7420};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7390} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7363} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7272};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7203} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7590} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7559};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7145} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6994};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[11], float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7077} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7316} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7702};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6920};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7321);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6976} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6948} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6860};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7543} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7514} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7047};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7064} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7096} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7449};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7378} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6881};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6317 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6421} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6491} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6354};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6288} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6222};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6197} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6232} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6231};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26499} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26473} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26504};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26452} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26468};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8946, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8770} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9035};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009} = {1'B0, N13666} + {1'B0, N13668} + {1'B0, N13670};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918;
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[11], float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26449} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26496} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26455};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100} = {1'B0, N13693} + {1'B0, N13695} + {1'B0, N13697};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7450} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7418} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7509};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7351} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7267} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6851};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3456 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3412 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7627);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7358} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7387};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7037} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7007} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6886};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7012} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7430} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7396};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6901} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6931} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7284};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6372);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6244 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6412} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6275};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7050);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7034} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6972};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7501} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7577};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[7], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7659} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7234} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7623};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3503 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7004} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7094} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7065};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[6], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[5]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6999} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7080} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7466};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[6] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[5] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[5] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[5]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8760};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8671};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26461} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26444};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6509 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6434 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6227);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6298);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6334} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6268};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6207} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6433};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6466} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6243} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6390};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7483} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6949} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7334};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26458} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26439};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26474} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26464} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26490};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8607, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26481} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26436} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26486};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9283 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[4] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6359 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6492);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[4]};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7354);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7506} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7476};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3603 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7558} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7534} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7417};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[5], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7612} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7305} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7115};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[5]};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9088};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[7]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8999};
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[8]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[8]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8901};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7663);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N3142 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3], float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7148};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2] & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655 = ((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7350 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N6885) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7310) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N7085;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[2] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8655 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8931) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8756);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9248) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9210)) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[3]) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[3]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[4] | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9024);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8926 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8822) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8668);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9158) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8636)) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8593) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8934));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9252 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8824);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9006 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8734) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8562);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9059) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8617)) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9162) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8738));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8892 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8639) | (!(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9061 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8642)));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8797 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9285;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8579 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9165) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8971)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8795);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9130 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8711 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9203);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762 = !((N13682 & N13680) | N13678);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868 = N13673 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708 = N13673 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9100;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8868) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8762)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8708);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9260 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9009);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8836 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9199) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9034);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9176 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8918;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8930) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8769)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8606);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9072 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8807);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26553 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26548) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8944);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26556 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26562;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26561) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26563)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26565);
assign {float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850} = {1'B0, N13440} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26200} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26247};
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9211 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8850);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9019 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8667);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9288;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8820 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9223);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8638 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9032);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9202;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9197 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8833);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9007 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8653);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13738;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8805 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9209);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8619 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9017);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9010;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8818 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9182);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8634 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8991);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8790 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9193);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8600 | N13310);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8983)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8806);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8889 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8802 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9168);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8613 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8978);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268 = !((N12784 & N13191) | N13189);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9180 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8773);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8988 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8581);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9185 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268) & (!N14065)) | (!N13085);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26158 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26147);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8597 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8963);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9164 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8764);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8976 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8567);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8604 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8969)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8793);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993 & N13012) | N13010);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9030)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8861);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26710) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26703);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[39] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842 & N12502) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842) & N12500);
assign x[22] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[39]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8566 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9161));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8679 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9242 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8601;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9080 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8939 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9258;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[38] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842 & N12495) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842) & N12493);
assign x[21] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[38]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8998 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8826));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8752 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8584 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9183) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[37] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842 & N12488) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842) & N12486);
assign x[20] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[37]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9090 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8933));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8736 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8688)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9015 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8665;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8846 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8992 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8721;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8778);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9092);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8632);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8727;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9217 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8859) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9122);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8598 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8568) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8828);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8622 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9156) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8993);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26140);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[35] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263 & N12481) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263) & N12479);
assign x[18] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[35]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8759 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8596));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9057 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9265 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9112;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9108 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8691 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8897;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[34] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263 & N12474) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263) & N12472);
assign x[17] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[34]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9189 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9023));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8774 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8616 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8719) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[33] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263 & N12467) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9263) & N12465);
assign x[16] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[33]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8857 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8698));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26737 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26170;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26165 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26143 | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26156));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26168) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26151 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[32] = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149 & N12547) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26149) & N12549));
assign x[15] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[32]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8746 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9273 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9120));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877 = !N14033;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9086 | N13026);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8877)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040 = (!N14061) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9174;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879 = N14061 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9237;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9220);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9154;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9053) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9125)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8964);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8743) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8570);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[31] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8879) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9040);
assign x[14] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[31]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9198 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8960 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8783));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8695 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292 = (!N12762) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8867;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140 = N12762 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9268;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[30] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9140) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9292);
assign x[13] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[30]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9008 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8630 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9214));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803 = (!N12772) ^ N12782;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651 = (!N12772) ^ N12784;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[29] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8651) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8803);
assign x[12] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[29]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259 = !(N12782 & (!N12784));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[28] = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9259 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8951;
assign x[11] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[28]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8724 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9299));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8696 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9065)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8929;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9247 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9011;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8741;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8894);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004 = ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8730) & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8789)) | (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8635);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612 = !((float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9167 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903) | float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9004);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[27] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8911) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9068);
assign x[10] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[27]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9150 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8986));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9071 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8625;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8956 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8917;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[26] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9170) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8572);
assign x[9] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[26]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8811 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8661));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9284) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[25] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8677) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8831);
assign x[8] = !((N14307 & N14309) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[25]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9239 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9075));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[24] = float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8796 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8612;
assign x[7] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[24]));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8922 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8750));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9060) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[23] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9096) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8940);
assign x[6] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[23] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8578 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9179));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[22] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8674) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8563;
assign x[5] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[22] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9013 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8839));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8823;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[21] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8602) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9195);
assign x[4] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[21] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8686 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9262));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[20] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9094) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9087;
assign x[3] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[20] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9103 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8949));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8592;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9064;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643 = !float_div_cynw_cm_float_rcp_E8_M23_0_inst_N13851;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[19] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8863) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8705);
assign x[2] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[19] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8772 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8610));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[18] = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8854) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8643;
assign x[1] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[18] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9206 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9038));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8715) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126 = (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8873) ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9117;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[17] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9126) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8903) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8967);
assign x[0] = !((N14309 & N14307) | (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[17] & N14305));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26692 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8670 & (!float_div_cynw_cm_float_rcp_E8_M23_0_inst_N9251));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698 = N12569 ^ float_div_cynw_cm_float_rcp_E8_M23_0_inst_N8842;
assign x[19] = !((N14309 & N14307) | (N14305 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_N26698));
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38 = float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38 | float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__33);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[30] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[7]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[29] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[6]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[28] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[5]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[27] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[4]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[26] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[3]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[25] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[2]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[24] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[1]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[23] = (float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__22[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[31] = !(float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__29 | (!a_sign));
reg x_reg_23__I2481_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__I2481_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[23];
	end
assign x[23] = x_reg_23__I2481_QOUT;
reg x_reg_24__I2482_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__I2482_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[24];
	end
assign x[24] = x_reg_24__I2482_QOUT;
reg x_reg_25__I2483_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__I2483_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[25];
	end
assign x[25] = x_reg_25__I2483_QOUT;
reg x_reg_26__I2484_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__I2484_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[26];
	end
assign x[26] = x_reg_26__I2484_QOUT;
reg x_reg_27__I2485_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__I2485_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[27];
	end
assign x[27] = x_reg_27__I2485_QOUT;
reg x_reg_28__I2486_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I2486_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[28];
	end
assign x[28] = x_reg_28__I2486_QOUT;
reg x_reg_29__I2487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__I2487_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[29];
	end
assign x[29] = x_reg_29__I2487_QOUT;
reg x_reg_30__I2488_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I2488_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[30];
	end
assign x[30] = x_reg_30__I2488_QOUT;
reg x_reg_31__I2489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2489_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[31];
	end
assign x[31] = x_reg_31__I2489_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[0] = x[0];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[1] = x[1];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[2] = x[2];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[3] = x[3];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[4] = x[4];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[5] = x[5];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[6] = x[6];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[7] = x[7];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[8] = x[8];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[9] = x[9];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[10] = x[10];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[11] = x[11];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[12] = x[12];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[13] = x[13];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__48[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[21] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[22] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[23] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__60[24] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_0_inst_inst_cellmath__64[36] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  s7LyQgDeqhk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



