/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:40:48 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755;
wire N4739,N4746,N4753,N4760,N4767,N4774,N4781 
	,N4788,N4795,N4802,N4809,N4816,N4823,N4830,N4837 
	,N4844,N4851,N4858,N4865,N4872,N4879,N4886,N4950 
	,N4952,N5188,N5201,N5203,N5227,N5229,N5313,N5318 
	,N5344,N5369,N5379,N5383,N5408,N5410,N5422,N5424 
	,N5431,N5433,N5440,N5449,N5458,N5476,N5858,N5910 
	,N5962,N6014,N6062,N6121,N6169,N6217,N6219,N6265 
	,N6313,N6361,N6409,N6452,N6568,N6577,N6582,N6584 
	,N6611,N6618,N6737,N6866,N6925,N6981,N7081,N7086 
	,N7114,N7118,N7234,N7242,N7248,N7250,N7256,N7258 
	,N7270,N7276,N7285,N7292,N7299,N7306,N7313,N7316 
	,N7327,N7337,N7339,N7345,N7355,N7357,N7363,N7373 
	,N7375,N7381,N7391,N7393,N7403,N7405,N7758,N8067 
	,N8068,N8069,N8233,N8240,N8244,N8246,N8249,N8264 
	,N8267,N8277,N8285,N8287,N8297,N8301,N8321,N8325 
	,N8329,N8330,N8334,N8339,N8347,N8353,N8355,N8356 
	,N8409,N8411,N8414,N8420,N8424,N8425,N8464,N8466 
	,N8471,N8474,N8489,N8493,N8494,N8500,N8503,N8504 
	,N8506,N8509,N8510,N8512,N8516,N8517,N8521,N8524 
	,N8550,N8553,N8556,N8557,N8559,N8562,N8563,N8570 
	,N8574,N8576,N8579,N8581,N8585,N8587,N8589,N8591 
	,N8593,N8596,N8598,N8601,N8603,N8606,N8642,N8643 
	,N8646,N8648,N8651,N8654,N8656,N8674,N8675,N8682 
	,N8684,N8685,N8687,N8690,N8693,N8704,N8711,N8718 
	,N8725,N8732,N8739,N8746;
reg x_reg_22__retimed_I4110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4110_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1];
	end
assign N7758 = x_reg_22__retimed_I4110_QOUT;
reg x_reg_0__retimed_I3953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3953_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669;
	end
assign N7405 = x_reg_0__retimed_I3953_QOUT;
reg x_reg_0__retimed_I3952_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3952_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15];
	end
assign N7403 = x_reg_0__retimed_I3952_QOUT;
reg x_reg_0__retimed_I3948_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3948_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670;
	end
assign N7393 = x_reg_0__retimed_I3948_QOUT;
reg x_reg_0__retimed_I3947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3947_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16];
	end
assign N7391 = x_reg_0__retimed_I3947_QOUT;
reg x_reg_0__retimed_I3943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3943_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588;
	end
assign N7381 = x_reg_0__retimed_I3943_QOUT;
reg x_reg_0__retimed_I3941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3941_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672;
	end
assign N7375 = x_reg_0__retimed_I3941_QOUT;
reg x_reg_0__retimed_I3940_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3940_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18];
	end
assign N7373 = x_reg_0__retimed_I3940_QOUT;
reg x_reg_0__retimed_I3936_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3936_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568;
	end
assign N7363 = x_reg_0__retimed_I3936_QOUT;
reg x_reg_0__retimed_I3934_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3934_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674;
	end
assign N7357 = x_reg_0__retimed_I3934_QOUT;
reg x_reg_0__retimed_I3933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3933_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20];
	end
assign N7355 = x_reg_0__retimed_I3933_QOUT;
reg x_reg_0__retimed_I3929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3929_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550;
	end
assign N7345 = x_reg_0__retimed_I3929_QOUT;
reg x_reg_0__retimed_I3927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3927_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676;
	end
assign N7339 = x_reg_0__retimed_I3927_QOUT;
reg x_reg_0__retimed_I3926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3926_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22];
	end
assign N7337 = x_reg_0__retimed_I3926_QOUT;
reg x_reg_0__retimed_I3922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3922_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533;
	end
assign N7327 = x_reg_0__retimed_I3922_QOUT;
reg x_reg_0__retimed_I3918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3918_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
	end
assign N7316 = x_reg_0__retimed_I3918_QOUT;
reg x_reg_0__retimed_I3917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3917_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539;
	end
assign N7313 = x_reg_0__retimed_I3917_QOUT;
reg x_reg_0__retimed_I3915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3915_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599;
	end
assign N7306 = x_reg_0__retimed_I3915_QOUT;
reg x_reg_0__retimed_I3913_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3913_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521;
	end
assign N7299 = x_reg_0__retimed_I3913_QOUT;
reg x_reg_0__retimed_I3911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3911_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581;
	end
assign N7292 = x_reg_0__retimed_I3911_QOUT;
reg x_reg_0__retimed_I3909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3909_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508;
	end
assign N7285 = x_reg_0__retimed_I3909_QOUT;
reg x_reg_0__retimed_I3906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3906_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24];
	end
assign N7276 = x_reg_0__retimed_I3906_QOUT;
reg x_reg_0__retimed_I3905_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3905_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562;
	end
assign N7270 = x_reg_0__retimed_I3905_QOUT;
reg x_reg_0__retimed_I3902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3902_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572;
	end
assign N7258 = x_reg_0__retimed_I3902_QOUT;
reg x_reg_0__retimed_I3901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3901_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593;
	end
assign N7256 = x_reg_0__retimed_I3901_QOUT;
reg x_reg_0__retimed_I3900_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3900_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630;
	end
assign N7250 = x_reg_0__retimed_I3900_QOUT;
reg x_reg_0__retimed_I3899_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3899_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589;
	end
assign N7248 = x_reg_0__retimed_I3899_QOUT;
reg x_reg_0__retimed_I3898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3898_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554;
	end
assign N7242 = x_reg_0__retimed_I3898_QOUT;
reg x_reg_0__retimed_I3896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3896_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614;
	end
assign N7234 = x_reg_0__retimed_I3896_QOUT;
reg x_reg_0__retimed_I3858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3858_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720;
	end
assign N7118 = x_reg_0__retimed_I3858_QOUT;
reg x_reg_0__retimed_I3856_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3856_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740;
	end
assign N7114 = x_reg_0__retimed_I3856_QOUT;
reg x_reg_0__retimed_I3844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3844_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789;
	end
assign N7086 = x_reg_0__retimed_I3844_QOUT;
reg x_reg_0__retimed_I3843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3843_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782;
	end
assign N7081 = x_reg_0__retimed_I3843_QOUT;
reg x_reg_0__retimed_I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3806_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751;
	end
assign N6981 = x_reg_0__retimed_I3806_QOUT;
reg x_reg_0__retimed_I3796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3796_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784;
	end
assign N6925 = x_reg_0__retimed_I3796_QOUT;
reg x_reg_0__retimed_I3785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3785_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733;
	end
assign N6866 = x_reg_0__retimed_I3785_QOUT;
reg x_reg_0__retimed_I3765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3765_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374;
	end
assign N6737 = x_reg_0__retimed_I3765_QOUT;
reg x_reg_0__retimed_I3736_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3736_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42;
	end
assign N6618 = x_reg_0__retimed_I3736_QOUT;
reg x_reg_0__retimed_I3733_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3733_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4;
	end
assign N6611 = x_reg_0__retimed_I3733_QOUT;
reg x_reg_0__retimed_I3723_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3723_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635;
	end
assign N6584 = x_reg_0__retimed_I3723_QOUT;
reg x_reg_0__retimed_I3722_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3722_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634;
	end
assign N6582 = x_reg_0__retimed_I3722_QOUT;
reg x_reg_0__retimed_I3720_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3720_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43;
	end
assign N6577 = x_reg_0__retimed_I3720_QOUT;
reg x_reg_0__retimed_I3716_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3716_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557;
	end
assign N6568 = x_reg_0__retimed_I3716_QOUT;
reg x_reg_6__retimed_I3680_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3680_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0];
	end
assign N6452 = x_reg_6__retimed_I3680_QOUT;
reg x_reg_7__retimed_I3663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3663_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1];
	end
assign N6409 = x_reg_7__retimed_I3663_QOUT;
reg x_reg_8__retimed_I3644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3644_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2];
	end
assign N6361 = x_reg_8__retimed_I3644_QOUT;
reg x_reg_9__retimed_I3625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3625_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3];
	end
assign N6313 = x_reg_9__retimed_I3625_QOUT;
reg x_reg_10__retimed_I3606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3606_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4];
	end
assign N6265 = x_reg_10__retimed_I3606_QOUT;
reg x_reg_11__retimed_I3588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3588_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13];
	end
assign N6219 = x_reg_11__retimed_I3588_QOUT;
reg x_reg_11__retimed_I3587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3587_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5];
	end
assign N6217 = x_reg_11__retimed_I3587_QOUT;
reg x_reg_12__retimed_I3568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3568_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6];
	end
assign N6169 = x_reg_12__retimed_I3568_QOUT;
reg x_reg_13__retimed_I3549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3549_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7];
	end
assign N6121 = x_reg_13__retimed_I3549_QOUT;
reg x_reg_14__retimed_I3529_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3529_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8];
	end
assign N6062 = x_reg_14__retimed_I3529_QOUT;
reg x_reg_15__retimed_I3510_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3510_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9];
	end
assign N6014 = x_reg_15__retimed_I3510_QOUT;
reg x_reg_16__retimed_I3489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3489_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10];
	end
assign N5962 = x_reg_16__retimed_I3489_QOUT;
reg x_reg_17__retimed_I3468_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3468_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11];
	end
assign N5910 = x_reg_17__retimed_I3468_QOUT;
reg x_reg_18__retimed_I3447_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3447_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12];
	end
assign N5858 = x_reg_18__retimed_I3447_QOUT;
reg x_reg_22__retimed_I3291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3291_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0];
	end
assign N5476 = x_reg_22__retimed_I3291_QOUT;
reg x_reg_22__retimed_I3285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3285_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605;
	end
assign N5458 = x_reg_22__retimed_I3285_QOUT;
reg x_reg_22__retimed_I3282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3282_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630;
	end
assign N5449 = x_reg_22__retimed_I3282_QOUT;
reg x_reg_22__retimed_I3279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3279_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600;
	end
assign N5440 = x_reg_22__retimed_I3279_QOUT;
reg x_reg_22__retimed_I3277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3277_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612;
	end
assign N5433 = x_reg_22__retimed_I3277_QOUT;
reg x_reg_22__retimed_I3276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3276_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622;
	end
assign N5431 = x_reg_22__retimed_I3276_QOUT;
reg x_reg_22__retimed_I3274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3274_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617;
	end
assign N5424 = x_reg_22__retimed_I3274_QOUT;
reg x_reg_22__retimed_I3273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3273_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5];
	end
assign N5422 = x_reg_22__retimed_I3273_QOUT;
reg x_reg_22__retimed_I3269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3269_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610;
	end
assign N5410 = x_reg_22__retimed_I3269_QOUT;
reg x_reg_22__retimed_I3268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3268_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6];
	end
assign N5408 = x_reg_22__retimed_I3268_QOUT;
reg x_reg_22__retimed_I3259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3259_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758;
	end
assign N5383 = x_reg_22__retimed_I3259_QOUT;
reg x_reg_22__retimed_I3258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3258_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134;
	end
assign N5379 = x_reg_22__retimed_I3258_QOUT;
reg x_reg_22__retimed_I3255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3255_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7];
	end
assign N5369 = x_reg_22__retimed_I3255_QOUT;
reg x_reg_22__retimed_I3244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3244_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189;
	end
assign N5344 = x_reg_22__retimed_I3244_QOUT;
reg x_reg_23__retimed_I3236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3236_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650;
	end
assign N5318 = x_reg_23__retimed_I3236_QOUT;
reg x_reg_7__retimed_I3234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3234_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790;
	end
assign N5313 = x_reg_7__retimed_I3234_QOUT;
reg x_reg_31__retimed_I3227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3227_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6;
	end
assign N5229 = x_reg_31__retimed_I3227_QOUT;
reg x_reg_31__retimed_I3226_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3226_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
	end
assign N5227 = x_reg_31__retimed_I3226_QOUT;
reg x_reg_23__retimed_I3218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3218_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12;
	end
assign N5203 = x_reg_23__retimed_I3218_QOUT;
reg x_reg_23__retimed_I3217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3217_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17;
	end
assign N5201 = x_reg_23__retimed_I3217_QOUT;
reg x_reg_22__retimed_I3215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
	end
assign N5188 = x_reg_22__retimed_I3215_QOUT;
reg x_reg_31__retimed_I3120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3120_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001;
	end
assign N4952 = x_reg_31__retimed_I3120_QOUT;
reg x_reg_31__retimed_I3119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3119_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010;
	end
assign N4950 = x_reg_31__retimed_I3119_QOUT;
reg x_reg_0__retimed_I3092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3092_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0];
	end
assign N4886 = x_reg_0__retimed_I3092_QOUT;
reg x_reg_1__retimed_I3089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3089_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1];
	end
assign N4879 = x_reg_1__retimed_I3089_QOUT;
reg x_reg_2__retimed_I3086_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3086_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2];
	end
assign N4872 = x_reg_2__retimed_I3086_QOUT;
reg x_reg_3__retimed_I3083_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3083_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3];
	end
assign N4865 = x_reg_3__retimed_I3083_QOUT;
reg x_reg_4__retimed_I3080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3080_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4];
	end
assign N4858 = x_reg_4__retimed_I3080_QOUT;
reg x_reg_5__retimed_I3077_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3077_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5];
	end
assign N4851 = x_reg_5__retimed_I3077_QOUT;
reg x_reg_6__retimed_I3074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3074_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6];
	end
assign N4844 = x_reg_6__retimed_I3074_QOUT;
reg x_reg_7__retimed_I3071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7];
	end
assign N4837 = x_reg_7__retimed_I3071_QOUT;
reg x_reg_8__retimed_I3068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8];
	end
assign N4830 = x_reg_8__retimed_I3068_QOUT;
reg x_reg_9__retimed_I3065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3065_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9];
	end
assign N4823 = x_reg_9__retimed_I3065_QOUT;
reg x_reg_10__retimed_I3062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3062_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10];
	end
assign N4816 = x_reg_10__retimed_I3062_QOUT;
reg x_reg_11__retimed_I3059_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3059_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11];
	end
assign N4809 = x_reg_11__retimed_I3059_QOUT;
reg x_reg_12__retimed_I3056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3056_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12];
	end
assign N4802 = x_reg_12__retimed_I3056_QOUT;
reg x_reg_13__retimed_I3053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3053_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13];
	end
assign N4795 = x_reg_13__retimed_I3053_QOUT;
reg x_reg_14__retimed_I3050_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3050_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14];
	end
assign N4788 = x_reg_14__retimed_I3050_QOUT;
reg x_reg_15__retimed_I3047_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3047_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15];
	end
assign N4781 = x_reg_15__retimed_I3047_QOUT;
reg x_reg_16__retimed_I3044_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3044_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16];
	end
assign N4774 = x_reg_16__retimed_I3044_QOUT;
reg x_reg_17__retimed_I3041_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3041_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17];
	end
assign N4767 = x_reg_17__retimed_I3041_QOUT;
reg x_reg_18__retimed_I3038_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3038_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18];
	end
assign N4760 = x_reg_18__retimed_I3038_QOUT;
reg x_reg_19__retimed_I3035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3035_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19];
	end
assign N4753 = x_reg_19__retimed_I3035_QOUT;
reg x_reg_20__retimed_I3032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3032_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20];
	end
assign N4746 = x_reg_20__retimed_I3032_QOUT;
reg x_reg_21__retimed_I3029_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3029_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21];
	end
assign N4739 = x_reg_21__retimed_I3029_QOUT;
assign bdw_enable = !astall;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083 = !(a_exp[0] & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149 = !((a_exp[7] & a_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652 = !a_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653 | a_man[1]) | a_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106 = !(a_man[10] | a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125 = !(a_man[6] | a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114 = !(a_man[8] | a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134 = !(a_man[4] | a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168 = !(b_exp[0] & b_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157 = !((b_exp[7] & b_exp[6]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208 = !(((b_man[0] | b_man[1]) | b_man[2]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191 = !(b_man[10] | b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210 = !(b_man[6] | b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199 = !(b_man[8] | b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219 = !(b_man[4] | b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15 = !((((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25] = a_sign ^ b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062 = ((a_exp[0] | a_exp[7]) | a_exp[1]) | a_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075 = ((a_exp[5] | a_exp[3]) | a_exp[4]) | a_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040 = ((b_exp[0] | b_exp[7]) | b_exp[1]) | b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054 = ((b_exp[5] | b_exp[3]) | b_exp[4]) | b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563 = !b_exp[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562 = !b_exp[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561 = !b_exp[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560 = !b_exp[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559 = !b_exp[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558 = !b_exp[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557 = !b_exp[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556 = !b_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333 = a_exp[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]} = {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]} = {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]} = {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556} + {1'B0, a_exp[0]};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566} = {1'B0, a_exp[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364} + {1'B0, a_exp[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568} = {1'B0, a_exp[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569} = {1'B0, a_exp[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561} + {1'B0, a_exp[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562} + {1'B0, a_exp[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572} = {1'B0, a_exp[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638 = !a_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661 = b_man[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950 = !b_man[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633 = !(a_man[21] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642 = a_man[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 = !a_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 = !b_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386 = !a_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387 = !b_man[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369 = !b_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 = !a_man[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378 = !b_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384 = !a_man[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378 & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 = !b_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427 = !a_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428 = !b_man[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410 = !b_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 = !a_man[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419 = !b_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425 = !a_man[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419 & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287 = !b_man[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468 = !a_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469 = !b_man[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451 = !b_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 = !a_man[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461 = !b_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466 = !a_man[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461 & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 = !b_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 = !a_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 = !b_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346 = !a_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333 = !b_man[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351 = !b_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344 = !a_man[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975 = !b_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975 | a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980 = !a_man[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985 = !(b_man[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986 = !a_man[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973 = !(b_man[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981 = !b_man[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977 = !(a_man[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980 & b_man[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341);
assign N8704 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 | a_man[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317 = !((N8704 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323 & a_man[5]));
assign N8711 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 | b_man[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321 = !((N8711 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319 & b_man[6]));
assign N8718 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 | a_man[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471 = !((N8718 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310 & a_man[7]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455);
assign N8725 = a_man[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430 = !((N8725 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298) | (a_man[11] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414);
assign N8732 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 | a_man[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389 = !((N8732 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264 & a_man[15]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384)) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373);
assign N8739 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 | a_man[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494 = !((N8739 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241 & a_man[19]));
assign N8746 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 | b_man[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650 = !((N8746 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459 & b_man[20]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638 & b_man[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[20]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[19]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556 ^ a_exp[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & a_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46] = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083 = !(((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7])));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[8]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[13]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[12]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[11]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[10]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10] = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[9]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518) | (!(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593)) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586 = !((N7248 & N7250) | (!(N7403 | N7405)));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564 = ((!N7391) & (!N7393)) | ((!N7242) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564) ^ N7234;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586) ^ N7242;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] = (!N7250) ^ N7248;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14] = (!N7256) ^ N7258;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 = !(N6219 | N5858);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]);
assign N8244 = !(N7250 & N7248);
assign N8249 = !N7242;
assign N8246 = ((!N7405) & (!N7403)) | (!N8244);
assign N8240 = !N7391;
assign N8233 = !N7393;
assign N8648 = !N7373;
assign N8642 = !N7375;
assign N8656 = !(N8648 & N8642);
assign N8646 = !N7234;
assign N8643 = !((N8233 & N8240) | (N8249 & N8246));
assign N8651 = !(N8646 | N8643);
assign N8654 = !(N7381 | N8651);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512 = ((!N8654) & (!N7313)) | (!N8656);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544 = N8654;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21];
assign N8287 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512 & N7306) | N7363);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605 = N8287;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549 = ((!N7357) & (!N7355)) | ((!N7299) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549) ^ N7292;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605) ^ N7299;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512) ^ N7306;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544) ^ N7313;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549 & N7292) | N7345);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22] = (!N7285) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629;
assign N8285 = !N7337;
assign N8277 = !N7339;
assign N8297 = !(N8285 & N8277);
assign N8684 = !(N7299 | N8287);
assign N8687 = !(N7355 | N7357);
assign N8685 = !(N8687 | N8684);
assign N8690 = !N7292;
assign N8693 = !(N8690 | N8685);
assign N8682 = !N7285;
assign N8301 = ((!N8693) & (!N7345)) | (!N8682);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558 = !(N8297 & N8301);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695 & b_man[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695) & a_man[22]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558) ^ N7270;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49] = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558 & N7270) | N7327);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24] = (!N7276) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622;
assign N8675 = !(N7276 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622);
assign N8267 = !N7316;
assign N8264 = !N8675;
assign N8674 = !N8267;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25] = !((N8264 & N8674) | ((!N8264) & N8267));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743);
assign N8466 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780;
assign N8464 = !N7086;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 & N7081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788);
assign N8474 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730;
assign N8471 = !(N8474 | N8464);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158 = (N7086 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730) | N8466;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129 = !(N8471 | N8466);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802 & (!N7081));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780);
assign N8516 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1] = ((!N6925) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729)) | (!N8516);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 = !(((!N6866) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23] | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735 = N8264 ^ N8267;
assign N8330 = ((!N5858) & (!N7118)) | (!N7114);
assign N8339 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769);
assign N8347 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714) & (!N8330)) | (!N8339);
assign N8356 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799);
assign N8325 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24])) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735);
assign N8334 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743) & (!N8356)) | (!N8325);
assign N8329 = !N8334;
assign N8355 = !(N8347 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780);
assign N8321 = !(N6981 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729);
assign N8353 = !(N8355 & N8329);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135 = !(N8321 | N8353);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715));
assign N8067 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158;
assign N8068 = !N8067;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 & N6265;
assign N8069 = !N5383;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4] = !(N8069 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N5858);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135 & N6313;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N5910);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6062) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6452);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6121;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173 = N6361 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N5962);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102 = N6409 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6014);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6169;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6217;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6219);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031 = N6452 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6062);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6121);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6169);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6219) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6217);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N5858) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6265);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N5910) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6313);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N5962) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6361);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134 & N6014) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134) & N6409);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42) ^ fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630 = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 | (!a_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565 = b_sign & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585 = !rm[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547 = !rm[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585 & rm[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 = !(rm[1] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582 & b_sign) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582) & a_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2] = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1];
assign N8411 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059)) | (!N6737);
assign N8420 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567;
assign N8425 = !N6618;
assign N8424 = !((N8411 & N8425) | ((!N8411) & N8420));
assign N8414 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2] | N8424);
assign N8409 = !N6611;
assign N8512 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099);
assign N8489 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1] & N6577) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]) & N8512));
assign N8494 = !N6568;
assign N8510 = !(N8409 | N8414);
assign N8509 = !((N8494 | N6584) | N8510);
assign N8521 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567;
assign N8493 = !(N8521 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558));
assign N8506 = !N6618;
assign N8504 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558 | N8506);
assign N8517 = !N6584;
assign N8500 = !N6582;
assign N8524 = !(N8500 & N8517);
assign N8503 = ((!N8493) & (!N8504)) | (!N8524);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55 = ((!N8489) & (!N8509)) | (!N8503);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23], fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[4]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[3]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[6]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[7]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[5]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[1]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574 & b_exp[2]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574) & a_exp[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2] & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6];
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619};
assign {fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592};
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614 = !N7758;
assign {N8559, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]} = {1'B0, N5476} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]};
assign {N8581, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]} = {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023} + {1'B0, N8559};
assign {N8550, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]} = {1'B0, N5458} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079} + {1'B0, N8581};
assign {N8574, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]} = {1'B0, N5449} + {1'B0, N8068} + {1'B0, N8550};
assign {N8601, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]} = {1'B0, N5440} + {1'B0, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030} + {1'B0, N8574};
assign N8557 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5] = !(N5383 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755 | N5379);
assign {N8576, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]} = {1'B0, N5431} + {1'B0, N5433} + {1'B0, N8601};
assign {N8603, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]} = {1'B0, N5422} + {1'B0, N5424} + {1'B0, N8576};
assign {N8570, fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]} = {1'B0, N5408} + {1'B0, N5410} + {1'B0, N8603};
assign N8593 = !(N5369 | N8570);
assign N8606 = !(N5344 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]);
assign N8562 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62 | N8593);
assign N8563 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]);
assign N8579 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]);
assign N8596 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7];
assign N8598 = !(N8606 & N8562);
assign N8587 = !(N8563 & N8579);
assign N8556 = !N5369;
assign N8591 = !N8570;
assign N8585 = !((N8591 & N8556) | ((!N8591) & N5369));
assign N8553 = !(N8585 & N8596);
assign N8589 = !((N8587 | N8557) | N8553);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751 = !(N8598 | N8589);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 | (!N5188));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769 = !(rm[0] & rm[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7 = !(rm[2] | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653 = fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790 = !(((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70 = N5313 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 = !(N5188 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]));
assign x[22] = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860 & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[21]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[21]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]));
assign x[21] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4739);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[20]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[20]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]));
assign x[20] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4746);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[19]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[19]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]));
assign x[19] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4753);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[18]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[18]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]));
assign x[18] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4760);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[17]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[17]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]));
assign x[17] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4767);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[16]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[16]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]));
assign x[16] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4774);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[15]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[15]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]));
assign x[15] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4781);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[14]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[14]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]));
assign x[14] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4788);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[13]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[13]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]));
assign x[13] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4795);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[12]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[12]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]));
assign x[12] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4802);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[11]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[11]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]));
assign x[11] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4809);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[10]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[10]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]));
assign x[10] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4816);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[9]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[9]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]));
assign x[9] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4823);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[8]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[8]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]));
assign x[8] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4830);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[7]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[7]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]));
assign x[7] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4837);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[6]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[6]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]));
assign x[6] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4844);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[5]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[5]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]));
assign x[5] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4851);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[4]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[4]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]));
assign x[4] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4858);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[3]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[3]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]));
assign x[3] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4865);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[2]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[2]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]));
assign x[2] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4872);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_man[1]) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]));
assign x[1] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4879);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_man[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]));
assign x[0] = (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820 & N4886);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745 = ((N5203 | N5201) | N5188) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 = !fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751;
assign x[30] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]);
assign x[29] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]);
assign x[28] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]);
assign x[27] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]);
assign x[26] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]);
assign x[25] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]);
assign x[24] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650 = ((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651 = N5318 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0] = ((N5201 | N5203) | N5188) | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651;
assign x[23] = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748 = a_sign | b_sign;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6) | (a_sign & b_sign);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952 = !((fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13 & a_sign) | (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931 & b_sign));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710 = ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13) & (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18)) | (!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63) & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004 = (fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5] & N5229) | ((!fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]) & N5227);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010 = !(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63 | fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706);
assign x[31] = (N4950 & fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004) | ((!N4950) & N4952);
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[29] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLL4SQrcqx8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/


