/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:40:48 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755;
wire N4739,N4746,N4753,N4760,N4767,N4774,N4781 
	,N4788,N4795,N4802,N4809,N4816,N4823,N4830,N4837 
	,N4844,N4851,N4858,N4865,N4872,N4879,N4886,N4950 
	,N4952,N5188,N5201,N5203,N5227,N5229,N5313,N5318 
	,N5344,N5369,N5379,N5383,N5408,N5410,N5422,N5424 
	,N5431,N5433,N5440,N5449,N5458,N5476,N5858,N5910 
	,N5962,N6014,N6062,N6121,N6169,N6217,N6219,N6265 
	,N6313,N6361,N6409,N6452,N6568,N6577,N6582,N6584 
	,N6611,N6618,N6737,N6866,N6925,N6981,N7081,N7086 
	,N7114,N7118,N7234,N7242,N7248,N7250,N7256,N7258 
	,N7270,N7276,N7285,N7292,N7299,N7306,N7313,N7316 
	,N7327,N7337,N7339,N7345,N7355,N7357,N7363,N7373 
	,N7375,N7381,N7391,N7393,N7403,N7405,N7758,N8067 
	,N8068,N8069,N8233,N8240,N8244,N8246,N8249,N8264 
	,N8267,N8277,N8285,N8287,N8297,N8301,N8321,N8325 
	,N8329,N8330,N8334,N8339,N8347,N8353,N8355,N8356 
	,N8409,N8411,N8414,N8420,N8424,N8425,N8464,N8466 
	,N8471,N8474,N8489,N8493,N8494,N8500,N8503,N8504 
	,N8506,N8509,N8510,N8512,N8516,N8517,N8521,N8524 
	,N8550,N8553,N8556,N8557,N8559,N8562,N8563,N8570 
	,N8574,N8576,N8579,N8581,N8585,N8587,N8589,N8591 
	,N8593,N8596,N8598,N8601,N8603,N8606,N8642,N8643 
	,N8646,N8648,N8651,N8654,N8656,N8674,N8675,N8682 
	,N8684,N8685,N8687,N8690,N8693,N8704,N8711,N8718 
	,N8725,N8732,N8739,N8746;
reg x_reg_22__retimed_I4110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4110_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1];
	end
assign N7758 = x_reg_22__retimed_I4110_QOUT;
reg x_reg_0__retimed_I3953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3953_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669;
	end
assign N7405 = x_reg_0__retimed_I3953_QOUT;
reg x_reg_0__retimed_I3952_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3952_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15];
	end
assign N7403 = x_reg_0__retimed_I3952_QOUT;
reg x_reg_0__retimed_I3948_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3948_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670;
	end
assign N7393 = x_reg_0__retimed_I3948_QOUT;
reg x_reg_0__retimed_I3947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3947_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16];
	end
assign N7391 = x_reg_0__retimed_I3947_QOUT;
reg x_reg_0__retimed_I3943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3943_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588;
	end
assign N7381 = x_reg_0__retimed_I3943_QOUT;
reg x_reg_0__retimed_I3941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3941_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672;
	end
assign N7375 = x_reg_0__retimed_I3941_QOUT;
reg x_reg_0__retimed_I3940_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3940_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18];
	end
assign N7373 = x_reg_0__retimed_I3940_QOUT;
reg x_reg_0__retimed_I3936_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3936_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568;
	end
assign N7363 = x_reg_0__retimed_I3936_QOUT;
reg x_reg_0__retimed_I3934_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3934_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674;
	end
assign N7357 = x_reg_0__retimed_I3934_QOUT;
reg x_reg_0__retimed_I3933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3933_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20];
	end
assign N7355 = x_reg_0__retimed_I3933_QOUT;
reg x_reg_0__retimed_I3929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3929_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550;
	end
assign N7345 = x_reg_0__retimed_I3929_QOUT;
reg x_reg_0__retimed_I3927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3927_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676;
	end
assign N7339 = x_reg_0__retimed_I3927_QOUT;
reg x_reg_0__retimed_I3926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3926_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22];
	end
assign N7337 = x_reg_0__retimed_I3926_QOUT;
reg x_reg_0__retimed_I3922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3922_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533;
	end
assign N7327 = x_reg_0__retimed_I3922_QOUT;
reg x_reg_0__retimed_I3918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3918_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25];
	end
assign N7316 = x_reg_0__retimed_I3918_QOUT;
reg x_reg_0__retimed_I3917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3917_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539;
	end
assign N7313 = x_reg_0__retimed_I3917_QOUT;
reg x_reg_0__retimed_I3915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3915_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599;
	end
assign N7306 = x_reg_0__retimed_I3915_QOUT;
reg x_reg_0__retimed_I3913_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3913_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521;
	end
assign N7299 = x_reg_0__retimed_I3913_QOUT;
reg x_reg_0__retimed_I3911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3911_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581;
	end
assign N7292 = x_reg_0__retimed_I3911_QOUT;
reg x_reg_0__retimed_I3909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3909_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508;
	end
assign N7285 = x_reg_0__retimed_I3909_QOUT;
reg x_reg_0__retimed_I3906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3906_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24];
	end
assign N7276 = x_reg_0__retimed_I3906_QOUT;
reg x_reg_0__retimed_I3905_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3905_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562;
	end
assign N7270 = x_reg_0__retimed_I3905_QOUT;
reg x_reg_0__retimed_I3902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3902_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572;
	end
assign N7258 = x_reg_0__retimed_I3902_QOUT;
reg x_reg_0__retimed_I3901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3901_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593;
	end
assign N7256 = x_reg_0__retimed_I3901_QOUT;
reg x_reg_0__retimed_I3900_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3900_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630;
	end
assign N7250 = x_reg_0__retimed_I3900_QOUT;
reg x_reg_0__retimed_I3899_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3899_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589;
	end
assign N7248 = x_reg_0__retimed_I3899_QOUT;
reg x_reg_0__retimed_I3898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3898_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554;
	end
assign N7242 = x_reg_0__retimed_I3898_QOUT;
reg x_reg_0__retimed_I3896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3896_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614;
	end
assign N7234 = x_reg_0__retimed_I3896_QOUT;
reg x_reg_0__retimed_I3858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3858_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720;
	end
assign N7118 = x_reg_0__retimed_I3858_QOUT;
reg x_reg_0__retimed_I3856_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3856_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740;
	end
assign N7114 = x_reg_0__retimed_I3856_QOUT;
reg x_reg_0__retimed_I3844_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3844_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789;
	end
assign N7086 = x_reg_0__retimed_I3844_QOUT;
reg x_reg_0__retimed_I3843_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3843_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782;
	end
assign N7081 = x_reg_0__retimed_I3843_QOUT;
reg x_reg_0__retimed_I3806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3806_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751;
	end
assign N6981 = x_reg_0__retimed_I3806_QOUT;
reg x_reg_0__retimed_I3796_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3796_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784;
	end
assign N6925 = x_reg_0__retimed_I3796_QOUT;
reg x_reg_0__retimed_I3785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3785_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733;
	end
assign N6866 = x_reg_0__retimed_I3785_QOUT;
reg x_reg_0__retimed_I3765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3765_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374;
	end
assign N6737 = x_reg_0__retimed_I3765_QOUT;
reg x_reg_0__retimed_I3736_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3736_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42;
	end
assign N6618 = x_reg_0__retimed_I3736_QOUT;
reg x_reg_0__retimed_I3733_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3733_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4;
	end
assign N6611 = x_reg_0__retimed_I3733_QOUT;
reg x_reg_0__retimed_I3723_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3723_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635;
	end
assign N6584 = x_reg_0__retimed_I3723_QOUT;
reg x_reg_0__retimed_I3722_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3722_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634;
	end
assign N6582 = x_reg_0__retimed_I3722_QOUT;
reg x_reg_0__retimed_I3720_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3720_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43;
	end
assign N6577 = x_reg_0__retimed_I3720_QOUT;
reg x_reg_0__retimed_I3716_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3716_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557;
	end
assign N6568 = x_reg_0__retimed_I3716_QOUT;
reg x_reg_6__retimed_I3680_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3680_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0];
	end
assign N6452 = x_reg_6__retimed_I3680_QOUT;
reg x_reg_7__retimed_I3663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3663_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1];
	end
assign N6409 = x_reg_7__retimed_I3663_QOUT;
reg x_reg_8__retimed_I3644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3644_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2];
	end
assign N6361 = x_reg_8__retimed_I3644_QOUT;
reg x_reg_9__retimed_I3625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3625_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3];
	end
assign N6313 = x_reg_9__retimed_I3625_QOUT;
reg x_reg_10__retimed_I3606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3606_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4];
	end
assign N6265 = x_reg_10__retimed_I3606_QOUT;
reg x_reg_11__retimed_I3588_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3588_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13];
	end
assign N6219 = x_reg_11__retimed_I3588_QOUT;
reg x_reg_11__retimed_I3587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3587_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5];
	end
assign N6217 = x_reg_11__retimed_I3587_QOUT;
reg x_reg_12__retimed_I3568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3568_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6];
	end
assign N6169 = x_reg_12__retimed_I3568_QOUT;
reg x_reg_13__retimed_I3549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3549_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7];
	end
assign N6121 = x_reg_13__retimed_I3549_QOUT;
reg x_reg_14__retimed_I3529_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3529_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8];
	end
assign N6062 = x_reg_14__retimed_I3529_QOUT;
reg x_reg_15__retimed_I3510_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3510_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9];
	end
assign N6014 = x_reg_15__retimed_I3510_QOUT;
reg x_reg_16__retimed_I3489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3489_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10];
	end
assign N5962 = x_reg_16__retimed_I3489_QOUT;
reg x_reg_17__retimed_I3468_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3468_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11];
	end
assign N5910 = x_reg_17__retimed_I3468_QOUT;
reg x_reg_18__retimed_I3447_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3447_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12];
	end
assign N5858 = x_reg_18__retimed_I3447_QOUT;
reg x_reg_22__retimed_I3291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3291_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0];
	end
assign N5476 = x_reg_22__retimed_I3291_QOUT;
reg x_reg_22__retimed_I3285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3285_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605;
	end
assign N5458 = x_reg_22__retimed_I3285_QOUT;
reg x_reg_22__retimed_I3282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3282_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630;
	end
assign N5449 = x_reg_22__retimed_I3282_QOUT;
reg x_reg_22__retimed_I3279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3279_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600;
	end
assign N5440 = x_reg_22__retimed_I3279_QOUT;
reg x_reg_22__retimed_I3277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3277_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612;
	end
assign N5433 = x_reg_22__retimed_I3277_QOUT;
reg x_reg_22__retimed_I3276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3276_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622;
	end
assign N5431 = x_reg_22__retimed_I3276_QOUT;
reg x_reg_22__retimed_I3274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3274_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617;
	end
assign N5424 = x_reg_22__retimed_I3274_QOUT;
reg x_reg_22__retimed_I3273_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3273_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5];
	end
assign N5422 = x_reg_22__retimed_I3273_QOUT;
reg x_reg_22__retimed_I3269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3269_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610;
	end
assign N5410 = x_reg_22__retimed_I3269_QOUT;
reg x_reg_22__retimed_I3268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3268_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6];
	end
assign N5408 = x_reg_22__retimed_I3268_QOUT;
reg x_reg_22__retimed_I3259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3259_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758;
	end
assign N5383 = x_reg_22__retimed_I3259_QOUT;
reg x_reg_22__retimed_I3258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3258_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134;
	end
assign N5379 = x_reg_22__retimed_I3258_QOUT;
reg x_reg_22__retimed_I3255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3255_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7];
	end
assign N5369 = x_reg_22__retimed_I3255_QOUT;
reg x_reg_22__retimed_I3244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3244_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189;
	end
assign N5344 = x_reg_22__retimed_I3244_QOUT;
reg x_reg_23__retimed_I3236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3236_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650;
	end
assign N5318 = x_reg_23__retimed_I3236_QOUT;
reg x_reg_7__retimed_I3234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3234_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790;
	end
assign N5313 = x_reg_7__retimed_I3234_QOUT;
reg x_reg_31__retimed_I3227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3227_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6;
	end
assign N5229 = x_reg_31__retimed_I3227_QOUT;
reg x_reg_31__retimed_I3226_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3226_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48;
	end
assign N5227 = x_reg_31__retimed_I3226_QOUT;
reg x_reg_23__retimed_I3218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3218_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12;
	end
assign N5203 = x_reg_23__retimed_I3218_QOUT;
reg x_reg_23__retimed_I3217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3217_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17;
	end
assign N5201 = x_reg_23__retimed_I3217_QOUT;
reg x_reg_22__retimed_I3215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63;
	end
assign N5188 = x_reg_22__retimed_I3215_QOUT;
reg x_reg_31__retimed_I3120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3120_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001;
	end
assign N4952 = x_reg_31__retimed_I3120_QOUT;
reg x_reg_31__retimed_I3119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3119_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010;
	end
assign N4950 = x_reg_31__retimed_I3119_QOUT;
reg x_reg_0__retimed_I3092_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3092_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0];
	end
assign N4886 = x_reg_0__retimed_I3092_QOUT;
reg x_reg_1__retimed_I3089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3089_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1];
	end
assign N4879 = x_reg_1__retimed_I3089_QOUT;
reg x_reg_2__retimed_I3086_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3086_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2];
	end
assign N4872 = x_reg_2__retimed_I3086_QOUT;
reg x_reg_3__retimed_I3083_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3083_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3];
	end
assign N4865 = x_reg_3__retimed_I3083_QOUT;
reg x_reg_4__retimed_I3080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3080_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4];
	end
assign N4858 = x_reg_4__retimed_I3080_QOUT;
reg x_reg_5__retimed_I3077_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3077_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5];
	end
assign N4851 = x_reg_5__retimed_I3077_QOUT;
reg x_reg_6__retimed_I3074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3074_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6];
	end
assign N4844 = x_reg_6__retimed_I3074_QOUT;
reg x_reg_7__retimed_I3071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7];
	end
assign N4837 = x_reg_7__retimed_I3071_QOUT;
reg x_reg_8__retimed_I3068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8];
	end
assign N4830 = x_reg_8__retimed_I3068_QOUT;
reg x_reg_9__retimed_I3065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3065_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9];
	end
assign N4823 = x_reg_9__retimed_I3065_QOUT;
reg x_reg_10__retimed_I3062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3062_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10];
	end
assign N4816 = x_reg_10__retimed_I3062_QOUT;
reg x_reg_11__retimed_I3059_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3059_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11];
	end
assign N4809 = x_reg_11__retimed_I3059_QOUT;
reg x_reg_12__retimed_I3056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3056_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12];
	end
assign N4802 = x_reg_12__retimed_I3056_QOUT;
reg x_reg_13__retimed_I3053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3053_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13];
	end
assign N4795 = x_reg_13__retimed_I3053_QOUT;
reg x_reg_14__retimed_I3050_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3050_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14];
	end
assign N4788 = x_reg_14__retimed_I3050_QOUT;
reg x_reg_15__retimed_I3047_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3047_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15];
	end
assign N4781 = x_reg_15__retimed_I3047_QOUT;
reg x_reg_16__retimed_I3044_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3044_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16];
	end
assign N4774 = x_reg_16__retimed_I3044_QOUT;
reg x_reg_17__retimed_I3041_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3041_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17];
	end
assign N4767 = x_reg_17__retimed_I3041_QOUT;
reg x_reg_18__retimed_I3038_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3038_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18];
	end
assign N4760 = x_reg_18__retimed_I3038_QOUT;
reg x_reg_19__retimed_I3035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3035_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19];
	end
assign N4753 = x_reg_19__retimed_I3035_QOUT;
reg x_reg_20__retimed_I3032_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3032_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20];
	end
assign N4746 = x_reg_20__retimed_I3032_QOUT;
reg x_reg_21__retimed_I3029_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3029_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21];
	end
assign N4739 = x_reg_21__retimed_I3029_QOUT;
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I0 (.Y(bdw_enable), .A(astall));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149), .A(a_exp[7]), .B(a_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3085));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7149));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652), .A(a_man[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11652));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B(a_man[1]), .C(a_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3119));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134), .A(a_man[4]), .B(a_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3106), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3125), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3114), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3134));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3123), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3117), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3128), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3138));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157), .A(b_exp[7]), .B(b_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3170));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3168), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7157));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3204));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219), .A(b_man[4]), .B(b_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3210), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3199), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3219));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3208), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3202), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3213), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3223));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__10));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]));
OR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N547));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12062), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12075));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12040), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12054));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12189), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__12), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I46 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I47 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .A(b_exp[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I48 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .A(b_exp[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I49 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .A(b_exp[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I50 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .A(b_exp[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I51 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .A(b_exp[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I52 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558), .A(b_exp[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .A(b_exp[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .A(b_exp[0]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I56 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3333));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I57 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3327));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I58 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3348));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I59 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3319));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I60 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3343));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I61 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3362));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I62 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3337));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3330));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[7]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I66 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .B(a_exp[0]));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I67 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3321));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I68 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3364), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N558));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I69 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3338));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I70 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3358));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I71 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N561), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3331));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I72 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N562), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12635));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I73 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12652));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3627), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N572), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12518), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12499), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[1]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3617), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N566), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3604), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N569), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3597), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N568), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
OAI211X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3620), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N571), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3612), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N570), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[5]));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3655));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[4]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[2]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950), .A(b_man[21]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633), .A(a_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642), .A(a_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11950));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459), .A(a_man[20]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241), .A(b_man[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386), .A(a_man[18]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387), .A(b_man[18]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12387), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12386));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369), .A(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371), .A(a_man[17]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378), .A(b_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384), .A(a_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12369));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12378), .B(a_man[16]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264), .A(b_man[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427), .A(a_man[14]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428), .A(b_man[14]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12428), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12427));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410), .A(b_man[13]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412), .A(a_man[13]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419), .A(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425), .A(a_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12410));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12419), .B(a_man[12]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287), .A(b_man[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468), .A(a_man[10]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469), .A(b_man[10]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12469), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12468));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451), .A(b_man[9]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453), .A(a_man[9]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461), .A(b_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466), .A(a_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12451));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12461), .B(a_man[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310), .A(b_man[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319), .A(a_man[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323), .A(b_man[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346), .A(a_man[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333), .A(b_man[4]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351), .A(b_man[3]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344), .A(a_man[3]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12333), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12346));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975), .A(b_man[2]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11975), .B(a_man[2]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12344), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12351));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980), .A(a_man[1]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I156 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I157 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986), .A(a_man[2]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I158 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11986));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I159 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981), .A(b_man[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I160 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977), .A(a_man[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11981));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I161 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972), .A0(b_man[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11980), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11977));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I162 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11985), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11973), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11972));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I163 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12338), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12343));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12350), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12352));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12336), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12341));
OR2XL cmpoi_A_I4587 (.Y(N8704), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323), .B(a_man[5]));
AOI22XL cmpoi_A_I4588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12314), .A1(N8704), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12323), .B1(a_man[5]));
OR2XL cmpoi_A_I4589 (.Y(N8711), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319), .B(b_man[6]));
AOI22XL cmpoi_A_I4590 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12317), .A1(N8711), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12319), .B1(b_man[6]));
OR2XL cmpoi_A_I4591 (.Y(N8718), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310), .B(a_man[7]));
AOI22XL cmpoi_A_I4592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12321), .A1(N8718), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12310), .B1(a_man[7]));
AOI222X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12460), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12466), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12453), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12450), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12456), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12471));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12464), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12457), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12462));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12473), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12455));
OR2XL cmpoi_A_I4593 (.Y(N8725), .A(a_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287));
AOI22XL cmpoi_A_I4594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12298), .A1(N8725), .B0(a_man[11]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12287));
AOI222X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12420), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12425), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12412), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12409), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12415), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12430));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12423), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12416), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12421));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12432), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12414));
OR2XL cmpoi_A_I4595 (.Y(N8732), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264), .B(a_man[15]));
AOI22XL cmpoi_A_I4596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12275), .A1(N8732), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12264), .B1(a_man[15]));
AOI222X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12379), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12384), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12371), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12368), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12374), .C1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12389));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12382), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12375), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12380));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12391), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12373));
OR2XL cmpoi_A_I4597 (.Y(N8739), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241), .B(a_man[19]));
AOI22XL cmpoi_A_I4598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12252), .A1(N8739), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12241), .B1(a_man[19]));
OR2XL cmpoi_A_I4599 (.Y(N8746), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459), .B(b_man[20]));
AOI22XL cmpoi_A_I4600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3494), .A1(N8746), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3459), .B1(b_man[20]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12642), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12650));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12638), .B(b_man[22]));
AOI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12661), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12633), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12658), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12662));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12639));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N575));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004), .A(b_man[20]), .B(a_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016), .A(b_man[19]), .B(a_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N556), .B(a_exp[0]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12017), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12005), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3614));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12492));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .A(b_man[4]), .B(a_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .A(b_man[3]), .B(a_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .A(b_man[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12687));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12507));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .A(b_man[11]), .B(a_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .A(b_man[14]), .B(a_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .A(b_man[13]), .B(a_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[25]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12016));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12004));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[24]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3925), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3953), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3868), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3897), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3849), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3983), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3793), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3957), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3861), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3885), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3807), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3803), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3833));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3970));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3911));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3815), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[26]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3810), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3841), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3790), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3961), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3959));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3909), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3905), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3932));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3858));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3906), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[7]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3817));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3982));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3937), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3882), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3979));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3934), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[5]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4291), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4300));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12043), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12060), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12038));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3852), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3876), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3800), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3938), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3795), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3931));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3977));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3973), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3784));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3778), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3854), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3830), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3922));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3847));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3825), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12073), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12033), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12046), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12086));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12036), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12083));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3822), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3886), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3884));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3927), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3775), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3794), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3839));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3880), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3891));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3812), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3916));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3769));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3888));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3845));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3837), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3929));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3865));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3863));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[10]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4265), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4274));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12057), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12092), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12079));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3781), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3873));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3919), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3940), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3819), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3958));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3827), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3777), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3943));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3912), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3792));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3835), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3945), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3788));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3766), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3805));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[17]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3786));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3878));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3975));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[2]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4261), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4271));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3918), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3894), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3772), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3967));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3910));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3955), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4282));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4279), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4294));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12052), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12066), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12070));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12049), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12063));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12076), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12088));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12091));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3809));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3856), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[26]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[26]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__44), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3924), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3968), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[33]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12713));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3875), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[32]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3832));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3871), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[31]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12699));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3783));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3828), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[30]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[30]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3952));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3779), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[29]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3903), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3948), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[28]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[28]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3860), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3899), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[27]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[27]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[1]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N655), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4556), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4618));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[2]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N656));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[3]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N657), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[4]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N658));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[5]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N659), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[6]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N660));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N661), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[8]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N662));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3972), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3798), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[34]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4534), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4623));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4604), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4566));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4537), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4511));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4592), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4582));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4510), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4524));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4540), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4601));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4575), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4541));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4758), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3963), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3811), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[41]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4554), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3821), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3933), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[40]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3774), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[39]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12720));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3960), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[38]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[38]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3896), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3866), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[37]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12727));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I495 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3770), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[36]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[36]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3846), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3802));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[35]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12734));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[9]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N663), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4585), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4546));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[10]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N664));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[11]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N665), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[12]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N666));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]));
AOI2BB2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[13]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N667), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518));
OAI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4589), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4572), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4593), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[14]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N668));
CLKXOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4630), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[15]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3904));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4614), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]));
AOI2BB2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586), .A0N(N7403), .A1N(N7405), .B0(N7248), .B1(N7250));
OAI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564), .A0(N7391), .A1(N7393), .B0(N7242), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4564), .B(N7234));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4586), .B(N7242));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]));
XNOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .A(N7250), .B(N7248));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .A(N7256), .B(N7258));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4576), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4518));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4561), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4594));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802), .A(N6219), .B(N5858));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4529), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4530));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4631), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4609));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4782), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3974));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4521), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[20]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3877));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4599), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3785));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4539), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4588), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[17]));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4388 (.Y(N8244), .A(N7250), .B(N7248));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4390 (.Y(N8249), .A(N7242));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4391 (.Y(N8246), .A0(N7403), .A1(N7405), .B0(N8244));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4392 (.Y(N8240), .A(N7391));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4393 (.Y(N8233), .A(N7393));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4564 (.Y(N8648), .A(N7373));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4565 (.Y(N8642), .A(N7375));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4566 (.Y(N8656), .A(N8648), .B(N8642));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4567 (.Y(N8646), .A(N7234));
AOI22X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4568 (.Y(N8643), .A0(N8240), .A1(N8233), .B0(N8249), .B1(N8246));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4569 (.Y(N8651), .A(N8646), .B(N8643));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4570 (.Y(N8654), .A(N7381), .B(N8651));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .A0(N7313), .A1(N8654), .B0(N8656));
DLY1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4572 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544), .A(N8654));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[19]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3853));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4581), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4407 (.Y(N8287), .A0(N7306), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .B0(N7363));
BUFX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605), .A(N8287));
OAI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .A0(N7357), .A1(N7355), .B0(N7299), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .B(N7292));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4605), .B(N7299));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4512), .B(N7306));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4544), .B(N7313));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4550), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[21]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3944));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4508), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[22]));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629), .A0(N7292), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4549), .B0(N7345));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .A(N7285), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4629));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4417 (.Y(N8285), .A(N7337));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4418 (.Y(N8277), .A(N7339));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4419 (.Y(N8297), .A(N8285), .B(N8277));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4580 (.Y(N8684), .A(N7299), .B(N8287));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4581 (.Y(N8687), .A(N7355), .B(N7357));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4582 (.Y(N8685), .A(N8687), .B(N8684));
CLKINVX8 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4583 (.Y(N8690), .A(N7292));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4584 (.Y(N8693), .A(N8690), .B(N8685));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4585 (.Y(N8682), .A(N7285));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4586 (.Y(N8301), .A0(N7345), .A1(N8693), .B0(N8682));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .A(N8297), .B(N8301));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3695));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3823));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4562), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .B(N7270));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I579 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4205), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3816), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3914));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[49]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4328));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4533), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[23]));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I582 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622), .A0(N7270), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4558), .B0(N7327));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I583 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A(N7276), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4574 (.Y(N8675), .A(N7276), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4622));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4575 (.Y(N8267), .A(N7316));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4576 (.Y(N8264), .A(N8675));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4577 (.Y(N8674), .A(N8267));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]), .A(N8267), .B(N8674), .S0(N8264));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4504 (.Y(N8466), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4505 (.Y(N8464), .A(N7086));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802), .B(N7081));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4509 (.Y(N8474), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4510 (.Y(N8471), .A(N8474), .B(N8464));
AO21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .A1(N7086), .B0(N8466));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129), .A(N8471), .B(N8466));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4725), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4744));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4784), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4752), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4792), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4771));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728), .AN(N7081), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4802));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4738));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4717), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4728), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4747));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4745), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4766));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4795));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4773), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4756), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4775));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4730), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4514 (.Y(N8516), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4797));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .A1(N6925), .B0(N8516));
CLKINVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4733), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4760));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4788), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4724), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4761), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4781));
OA21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729), .A1(N6866), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4801));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I608 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I610 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I612 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4757), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4776));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I614 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4786), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4806));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4779), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4798), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4734));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4751), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4736), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4723));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4720), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4740), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[13]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I621 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I625 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]));
NOR2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735), .A(N8264), .B(N8267));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4430 (.Y(N8330), .A0(N7118), .A1(N5858), .B0(N7114));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4431 (.Y(N8339), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4748), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4769));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4432 (.Y(N8347), .A0(N8330), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4714), .B0(N8339));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4433 (.Y(N8356), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4777), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4799));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4434 (.Y(N8325), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4712), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4735));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4435 (.Y(N8334), .A0(N8356), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4743), .B0(N8325));
CLKINVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4436 (.Y(N8329), .A(N8334));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4437 (.Y(N8355), .A(N8347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4780));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4438 (.Y(N8321), .A(N6981), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4439 (.Y(N8353), .A(N8355), .B(N8329));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .A(N8321), .B(N8353));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11648));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11788));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4789), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4715), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4719));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4265 (.Y(N8067), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4266 (.Y(N8068), .A(N8067));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .B(N6265));
INVXL compensate_x_1_A_I4267 (.Y(N8069), .A(N5383));
NOR2XL compensate_x_1_A_I4268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4]), .A(N8069), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729));
CLKINVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I647 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7129));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I648 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047), .A(N5858), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I649 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5047), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I650 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135), .B(N6313));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176), .A(N5910), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5176), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135));
CLKINVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11650));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .A(N6452), .B(N6062), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5026), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(N6121));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I661 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[23]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5155), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5142), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5086), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173), .A(N6361), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139), .A(N5962), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102), .A(N6409), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7135));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105), .A(N6014), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5105), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(N6169));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I673 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5119), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134), .B(N6217));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084), .A(N6219), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5084), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5178), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
CLKINVX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5045), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5127), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5093), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5108), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5071), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5049), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031), .A(N6452), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5158));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068), .A(N6062), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5066), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5068), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5056), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5037), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5163), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I690 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I691 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5172), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I692 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034), .A(N6121), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I693 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5034), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I694 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5019), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I695 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5106), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I696 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5136), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I697 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160), .A(N6169), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I698 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5160), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I699 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5114), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I700 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5069), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I701 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5101), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124), .A(N6217), .B(N6219), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5124), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5043), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5036), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I706 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5065), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090), .A(N6265), .B(N5858), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5090), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5133), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5162), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053), .A(N6313), .B(N5910), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I713 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5053), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I714 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5063), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I715 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5126), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I716 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5157), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016), .A(N6361), .B(N5962), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5016), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5154), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5092), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5121), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146), .A(N6409), .B(N6014), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7134));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5146), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5083), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5054), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5087), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5111), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5175), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5017), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5050), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5040), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5104), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5148), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5179), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I735 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5130), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5033), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5113), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5143), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5060), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5123), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5076), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5109), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5151), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5052), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5042), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5072), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5080), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5145), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5167), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I750 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5038), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I751 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5173));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I752 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5074), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11789), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5131), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5102));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5166), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5098), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I758 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5128), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5031));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11649), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11651), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I761 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5062), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I762 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5094), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5022), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5116), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5025), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5057), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5153), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5020), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I768 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5117));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5149), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5081));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I771 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5077), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5138));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N626));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__30), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N628), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N627));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I779 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N630), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__39[25]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__32));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I782 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12695));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I783 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12595));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548), .AN(a_sign), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565), .A(b_sign), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .A(rm[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .A(rm[1]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .C(rm[0]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I789 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12548), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12565), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12547), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .C(rm[0]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12557), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12573), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5374), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__42), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__43));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12585), .B(rm[0]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5), .A(rm[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12741));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48), .A(a_sign), .B(b_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12582));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5169));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4455 (.Y(N8411), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12575), .B0(N6737));
CLKINVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4456 (.Y(N8420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4457 (.Y(N8425), .A(N6618));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4458 (.Y(N8424), .A(N8420), .B(N8425), .S0(N8411));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4459 (.Y(N8414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]), .B(N8424));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4460 (.Y(N8409), .A(N6611));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4519 (.Y(N8512), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5059), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5099));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4520 (.Y(N8489), .A(N8512), .B(N6577), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4521 (.Y(N8494), .A(N6568));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4522 (.Y(N8510), .A(N8409), .B(N8414));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4523 (.Y(N8509), .A(N8494), .B(N6584), .C(N8510));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4526 (.Y(N8521), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12567));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4527 (.Y(N8493), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558), .B(N8521));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4528 (.Y(N8506), .A(N6618));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4529 (.Y(N8504), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12558), .B(N8506));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4530 (.Y(N8517), .A(N6584));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4531 (.Y(N8500), .A(N6582));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4532 (.Y(N8524), .A(N8500), .B(N8517));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4533 (.Y(N8503), .A0(N8504), .A1(N8493), .B0(N8524));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55), .A0(N8509), .A1(N8489), .B0(N8503));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I810 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__55));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I811 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5477));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I812 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5466));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I813 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5456));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I814 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5449));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I815 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5438));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I816 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5429));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I817 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5421));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I818 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5482));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I819 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5474));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I820 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5464));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I821 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5454));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I822 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5446));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I823 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5436));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I824 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5428));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I825 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5418));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I826 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5480));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I827 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5473));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I828 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5461));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I829 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5452));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I830 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5445));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I831 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5434));
ADDHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I832 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5426));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12151), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[25]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N3367));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]), .A(a_exp[6]), .B(b_exp[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I840 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]), .A(a_exp[7]), .B(b_exp[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5584));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5583));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N574));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12134), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5580), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[6]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I851 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5605), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[2]));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I852 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5630), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5619));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I853 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5612), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5592));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5622), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__29[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614), .A(N7758));
ADDFXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4538 (.CO(N8559), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5135), .B(N5476), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[23]));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4539 (.CO(N8581), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5023), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5614), .CI(N8559));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4540 (.CO(N8550), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5079), .B(N5458), .CI(N8581));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4541 (.CO(N8574), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]), .A(N8068), .B(N5449), .CI(N8550));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4542 (.CO(N8601), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5030), .B(N5440), .CI(N8574));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4543 (.Y(N8557), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]), .A(N5383), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4729));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12755), .B(N5379));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4546 (.CO(N8576), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .A(N5433), .B(N5431), .CI(N8601));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4547 (.CO(N8603), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]), .A(N5424), .B(N5422), .CI(N8576));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4548 (.CO(N8570), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]), .A(N5410), .B(N5408), .CI(N8603));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4549 (.Y(N8593), .A(N5369), .B(N8570));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4550 (.Y(N8606), .A(N5344), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4551 (.Y(N8562), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .B(N8593));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4552 (.Y(N8563), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4553 (.Y(N8579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4554 (.Y(N8596), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4555 (.Y(N8598), .A(N8606), .B(N8562));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4556 (.Y(N8587), .A(N8563), .B(N8579));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4557 (.Y(N8556), .A(N5369));
CLKINVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4558 (.Y(N8591), .A(N8570));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4559 (.Y(N8585), .A(N5369), .B(N8556), .S0(N8591));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4560 (.Y(N8553), .A(N8585), .B(N8596));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4561 (.Y(N8589), .A(N8587), .B(N8557), .C(N8553));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I4562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751), .A(N8598), .B(N8589));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
CLKINVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
NOR2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .AN(N5188), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769), .A(rm[0]), .B(rm[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5769));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5354), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__5));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__7), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N652));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5790), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N653), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62), .B(N5313));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .A(N5188), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I885 (.Y(x[22]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5860));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[21]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[21]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[21]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I889 (.Y(x[21]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4739), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5817));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[20]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[20]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[20]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I892 (.Y(x[20]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4746), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5873));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I893 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[19]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I894 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[19]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I895 (.Y(x[19]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4753), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5831));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I896 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[18]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[18]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I897 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7139), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[18]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I898 (.Y(x[18]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4760), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5886));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I899 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[17]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I900 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I901 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[17]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I902 (.Y(x[17]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4767), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5844));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[16]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[16]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[16]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I905 (.Y(x[16]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4774), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5801));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I906 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[15]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[15]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I907 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[15]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I908 (.Y(x[15]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4781), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5856));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[14]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[14]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I911 (.Y(x[14]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4788), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5812));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[13]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7140), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I914 (.Y(x[13]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4795), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5868));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I915 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[12]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I916 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7138));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I918 (.Y(x[12]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4802), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5825));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[11]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[11]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I920 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I921 (.Y(x[11]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4809), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5881));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[10]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[10]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I923 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[10]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I924 (.Y(x[10]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4816), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5839));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I925 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[9]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[9]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I927 (.Y(x[9]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4823), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5796));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I928 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[8]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I929 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[8]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I930 (.Y(x[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4830), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5851));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[7]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I933 (.Y(x[7]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4837), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5808));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I935 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[6]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I936 (.Y(x[6]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4844), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5864));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I937 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I938 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[5]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I939 (.Y(x[5]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4851), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5821));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[4]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I942 (.Y(x[4]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4858), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5877));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[3]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I945 (.Y(x[3]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4865), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5834));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[2]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I948 (.Y(x[2]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4872), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5889));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(a_man[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[1]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I951 (.Y(x[1]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4879), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5847));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N11653), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_man[0]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5875), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N7143), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__57[0]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I954 (.Y(x[0]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5820), .A1N(N4886), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5804));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .A(N5203), .B(N5201), .C(N5188), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5751));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I957 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I958 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I959 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I960 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I961 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I962 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I963 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5745), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I964 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__4), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N634), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N635));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651), .A(N5318), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__62));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]), .A(N5201), .B(N5203), .C(N5188), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I967 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5733));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I968 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748), .A(a_sign), .B(b_sign));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N12748), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__16), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N645));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952), .A0(a_sign), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4931), .B1(b_sign));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__18), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N4952));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5001), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I974 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004), .A(N5227), .B(N5229), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5010), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_3_I976 (.Y(x[31]), .A(N4952), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_N5004), .S0(N4950));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[29] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__33[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__50[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_2_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  uLn1TAHaqhE= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/


