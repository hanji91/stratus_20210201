/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:06:59 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
wire N11500,N11504,N11506,N11667,N11672,N11677,N11682 
	,N11687,N11692,N11697,N11702,N11707,N11712,N11717,N11722 
	,N11788,N11798,N11806,N11814,N11822,N11830,N11838,N11846 
	,N11854,N11862,N11886,N11937,N11941,N11966,N12003,N12007 
	,N12042,N12044,N12077,N12085,N12087,N12089,N12122,N12130 
	,N12132,N12167,N12169,N12175,N12177,N12183,N12218,N12220 
	,N12238,N12240,N12242,N12277,N12279,N12285,N12289,N12293 
	,N12295,N12297,N12325,N12327,N12363,N12365,N12383,N12413 
	,N12415,N12421,N12423,N12429,N12435,N12443,N12445,N12447 
	,N12480,N12482,N12488,N12490,N12492,N12496,N12498,N12500 
	,N12504,N12506,N12508,N12512,N12514,N12516,N12529,N12542 
	,N12544,N12550,N12552,N12554,N12560,N12562,N12564,N12567 
	,N12578,N12580,N12582,N12585,N12587,N12589,N12591,N12605 
	,N12607,N12609,N12613,N12618,N12625,N12627,N13149,N13150 
	,N13151,N13152,N13153,N13154,N13155,N13156,N13164,N13166 
	,N13167,N13170,N13172,N13174,N13178,N13180,N13181,N13182 
	,N13202,N13204,N13205,N13209,N13212,N13215,N13229,N13232 
	,N13234,N13236,N13238,N13241,N13242,N13246,N13248,N13250 
	,N13251,N13254,N13256,N13259,N13263,N13264,N13266,N13267 
	,N13268,N13269,N13271,N13273,N13274,N13277,N13279,N13281 
	,N13318,N13319,N13322,N13326,N13329,N13330,N13337,N13353 
	,N13354,N13356,N13358,N13359,N13360,N13362,N13364,N13366 
	,N13368,N13370,N13371,N13373,N13376,N13378,N13380,N13382 
	,N13385,N13389,N13391,N13392,N13395,N13400,N13436,N13440 
	,N13443,N13445,N13447,N13450,N13452,N13455,N13457,N13459 
	,N13460,N13461,N13463,N13464,N13466,N13468,N13470,N13472 
	,N13474,N13476,N13478,N13479,N13482,N13484,N13486,N13518 
	,N13521,N13530,N13542,N13543,N13546,N13548,N13550,N13551 
	,N13553,N13556,N13557,N13562,N13564,N13566,N13568,N13570 
	,N13571,N13573,N13575,N13577,N13579,N13581,N13583,N13586 
	,N13588,N13590,N13591,N13626,N13628,N13630,N13632,N13634 
	,N13636,N13639,N13642,N13645,N13647,N13649,N13650,N13651 
	,N13653,N13655,N13659,N13661,N13663,N13665,N13667,N13668 
	,N13671;
reg x_reg_22__retimed_I7284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7284_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14];
	end
assign N12627 = x_reg_22__retimed_I7284_QOUT;
reg x_reg_22__retimed_I7283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7283_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13];
	end
assign N12625 = x_reg_22__retimed_I7283_QOUT;
reg x_reg_22__retimed_I7278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648;
	end
assign N12609 = x_reg_22__retimed_I7278_QOUT;
reg x_reg_22__retimed_I7277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7277_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832;
	end
assign N12607 = x_reg_22__retimed_I7277_QOUT;
reg x_reg_22__retimed_I7276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7276_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11];
	end
assign N12605 = x_reg_22__retimed_I7276_QOUT;
reg x_reg_22__retimed_I7272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7272_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564;
	end
assign N12591 = x_reg_22__retimed_I7272_QOUT;
reg x_reg_22__retimed_I7271_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7271_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570;
	end
assign N12589 = x_reg_22__retimed_I7271_QOUT;
reg x_reg_22__retimed_I7270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7270_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919;
	end
assign N12587 = x_reg_22__retimed_I7270_QOUT;
reg x_reg_22__retimed_I7269_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7269_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800;
	end
assign N12585 = x_reg_22__retimed_I7269_QOUT;
reg x_reg_22__retimed_I7268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7268_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13];
	end
assign N12582 = x_reg_22__retimed_I7268_QOUT;
reg x_reg_22__retimed_I7267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7267_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13];
	end
assign N12580 = x_reg_22__retimed_I7267_QOUT;
reg x_reg_22__retimed_I7266_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7266_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13];
	end
assign N12578 = x_reg_22__retimed_I7266_QOUT;
reg x_reg_22__retimed_I7262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7262_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703;
	end
assign N12567 = x_reg_22__retimed_I7262_QOUT;
reg x_reg_22__retimed_I7261_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7261_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12];
	end
assign N12564 = x_reg_22__retimed_I7261_QOUT;
reg x_reg_22__retimed_I7260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7260_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550;
	end
assign N12562 = x_reg_22__retimed_I7260_QOUT;
reg x_reg_22__retimed_I7259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7259_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622;
	end
assign N12560 = x_reg_22__retimed_I7259_QOUT;
reg x_reg_22__retimed_I7258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7258_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359;
	end
assign N12554 = x_reg_22__retimed_I7258_QOUT;
reg x_reg_22__retimed_I7257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7257_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265;
	end
assign N12552 = x_reg_22__retimed_I7257_QOUT;
reg x_reg_22__retimed_I7256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7256_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209;
	end
assign N12550 = x_reg_22__retimed_I7256_QOUT;
reg x_reg_22__retimed_I7254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7254_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14];
	end
assign N12544 = x_reg_22__retimed_I7254_QOUT;
reg x_reg_22__retimed_I7253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14];
	end
assign N12542 = x_reg_22__retimed_I7253_QOUT;
reg x_reg_22__retimed_I7248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7248_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024;
	end
assign N12529 = x_reg_22__retimed_I7248_QOUT;
reg x_reg_22__retimed_I7244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7244_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295;
	end
assign N12516 = x_reg_22__retimed_I7244_QOUT;
reg x_reg_22__retimed_I7243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7243_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283;
	end
assign N12514 = x_reg_22__retimed_I7243_QOUT;
reg x_reg_22__retimed_I7242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7242_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149;
	end
assign N12512 = x_reg_22__retimed_I7242_QOUT;
reg x_reg_22__retimed_I7241_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7241_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275;
	end
assign N12508 = x_reg_22__retimed_I7241_QOUT;
reg x_reg_22__retimed_I7240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7240_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075;
	end
assign N12506 = x_reg_22__retimed_I7240_QOUT;
reg x_reg_22__retimed_I7239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7239_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128;
	end
assign N12504 = x_reg_22__retimed_I7239_QOUT;
reg x_reg_22__retimed_I7238_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7238_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351;
	end
assign N12500 = x_reg_22__retimed_I7238_QOUT;
reg x_reg_22__retimed_I7237_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7237_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257;
	end
assign N12498 = x_reg_22__retimed_I7237_QOUT;
reg x_reg_22__retimed_I7236_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7236_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203;
	end
assign N12496 = x_reg_22__retimed_I7236_QOUT;
reg x_reg_22__retimed_I7235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7235_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184;
	end
assign N12492 = x_reg_22__retimed_I7235_QOUT;
reg x_reg_22__retimed_I7234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7234_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378;
	end
assign N12490 = x_reg_22__retimed_I7234_QOUT;
reg x_reg_22__retimed_I7233_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7233_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092;
	end
assign N12488 = x_reg_22__retimed_I7233_QOUT;
reg x_reg_22__retimed_I7231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7231_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15];
	end
assign N12482 = x_reg_22__retimed_I7231_QOUT;
reg x_reg_22__retimed_I7230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7230_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487;
	end
assign N12480 = x_reg_22__retimed_I7230_QOUT;
reg x_reg_22__retimed_I7218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7218_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167;
	end
assign N12447 = x_reg_22__retimed_I7218_QOUT;
reg x_reg_22__retimed_I7217_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7217_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358;
	end
assign N12445 = x_reg_22__retimed_I7217_QOUT;
reg x_reg_22__retimed_I7216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7216_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343;
	end
assign N12443 = x_reg_22__retimed_I7216_QOUT;
reg x_reg_22__retimed_I7213_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7213_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090;
	end
assign N12435 = x_reg_22__retimed_I7213_QOUT;
reg x_reg_22__retimed_I7211_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7211_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16];
	end
assign N12429 = x_reg_22__retimed_I7211_QOUT;
reg x_reg_22__retimed_I7209_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7209_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083;
	end
assign N12423 = x_reg_22__retimed_I7209_QOUT;
reg x_reg_22__retimed_I7208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7208_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223;
	end
assign N12421 = x_reg_22__retimed_I7208_QOUT;
reg x_reg_22__retimed_I7206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7206_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757;
	end
assign N12415 = x_reg_22__retimed_I7206_QOUT;
reg x_reg_22__retimed_I7205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7205_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618;
	end
assign N12413 = x_reg_22__retimed_I7205_QOUT;
reg x_reg_22__retimed_I7194_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7194_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155;
	end
assign N12383 = x_reg_22__retimed_I7194_QOUT;
reg x_reg_22__retimed_I7188_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7188_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945;
	end
assign N12365 = x_reg_22__retimed_I7188_QOUT;
reg x_reg_22__retimed_I7187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7187_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890;
	end
assign N12363 = x_reg_22__retimed_I7187_QOUT;
reg x_reg_22__retimed_I7174_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7174_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864;
	end
assign N12327 = x_reg_22__retimed_I7174_QOUT;
reg x_reg_22__retimed_I7173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7173_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457;
	end
assign N12325 = x_reg_22__retimed_I7173_QOUT;
reg x_reg_22__retimed_I7163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7163_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288;
	end
assign N12297 = x_reg_22__retimed_I7163_QOUT;
reg x_reg_22__retimed_I7162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7162_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317;
	end
assign N12295 = x_reg_22__retimed_I7162_QOUT;
reg x_reg_22__retimed_I7161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7161_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143;
	end
assign N12293 = x_reg_22__retimed_I7161_QOUT;
reg x_reg_22__retimed_I7160_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7160_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213;
	end
assign N12289 = x_reg_22__retimed_I7160_QOUT;
reg x_reg_22__retimed_I7158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7158_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228;
	end
assign N12285 = x_reg_22__retimed_I7158_QOUT;
reg x_reg_22__retimed_I7156_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7156_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787;
	end
assign N12279 = x_reg_22__retimed_I7156_QOUT;
reg x_reg_22__retimed_I7155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7155_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001;
	end
assign N12277 = x_reg_22__retimed_I7155_QOUT;
reg x_reg_22__retimed_I7143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7143_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392;
	end
assign N12242 = x_reg_22__retimed_I7143_QOUT;
reg x_reg_22__retimed_I7142_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7142_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272;
	end
assign N12240 = x_reg_22__retimed_I7142_QOUT;
reg x_reg_22__retimed_I7141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7141_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244;
	end
assign N12238 = x_reg_22__retimed_I7141_QOUT;
reg x_reg_22__retimed_I7135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7135_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709;
	end
assign N12220 = x_reg_22__retimed_I7135_QOUT;
reg x_reg_22__retimed_I7134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7134_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924;
	end
assign N12218 = x_reg_22__retimed_I7134_QOUT;
reg x_reg_22__retimed_I7122_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7122_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22];
	end
assign N12183 = x_reg_22__retimed_I7122_QOUT;
reg x_reg_22__retimed_I7120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7120_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22];
	end
assign N12177 = x_reg_22__retimed_I7120_QOUT;
reg x_reg_22__retimed_I7119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7119_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484;
	end
assign N12175 = x_reg_22__retimed_I7119_QOUT;
reg x_reg_22__retimed_I7117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7117_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627;
	end
assign N12169 = x_reg_22__retimed_I7117_QOUT;
reg x_reg_22__retimed_I7116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7116_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838;
	end
assign N12167 = x_reg_22__retimed_I7116_QOUT;
reg x_reg_22__retimed_I7104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7104_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23];
	end
assign N12132 = x_reg_22__retimed_I7104_QOUT;
reg x_reg_22__retimed_I7103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7103_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485;
	end
assign N12130 = x_reg_22__retimed_I7103_QOUT;
reg x_reg_22__retimed_I7100_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7100_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767;
	end
assign N12122 = x_reg_22__retimed_I7100_QOUT;
reg x_reg_22__retimed_I7089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7089_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24];
	end
assign N12089 = x_reg_22__retimed_I7089_QOUT;
reg x_reg_22__retimed_I7088_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7088_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24];
	end
assign N12087 = x_reg_22__retimed_I7088_QOUT;
reg x_reg_22__retimed_I7087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7087_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486;
	end
assign N12085 = x_reg_22__retimed_I7087_QOUT;
reg x_reg_22__retimed_I7084_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7084_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741;
	end
assign N12077 = x_reg_22__retimed_I7084_QOUT;
reg x_reg_22__retimed_I7073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7073_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874;
	end
assign N12044 = x_reg_22__retimed_I7073_QOUT;
reg x_reg_22__retimed_I7072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7072_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659;
	end
assign N12042 = x_reg_22__retimed_I7072_QOUT;
reg x_reg_22__retimed_I7060_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7060_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795;
	end
assign N12007 = x_reg_22__retimed_I7060_QOUT;
reg x_reg_22__retimed_I7058_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7058_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487;
	end
assign N12003 = x_reg_22__retimed_I7058_QOUT;
reg x_reg_22__retimed_I7045_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7045_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585;
	end
assign N11966 = x_reg_22__retimed_I7045_QOUT;
reg x_reg_22__retimed_I7037_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7037_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982;
	end
assign N11941 = x_reg_22__retimed_I7037_QOUT;
reg x_reg_22__retimed_I7035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7035_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719;
	end
assign N11937 = x_reg_22__retimed_I7035_QOUT;
reg x_reg_22__retimed_I7017_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7017_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638;
	end
assign N11886 = x_reg_22__retimed_I7017_QOUT;
reg x_reg_22__retimed_I7008_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7008_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976;
	end
assign N11862 = x_reg_22__retimed_I7008_QOUT;
reg x_reg_22__retimed_I7005_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7005_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683;
	end
assign N11854 = x_reg_22__retimed_I7005_QOUT;
reg x_reg_22__retimed_I7002_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I7002_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009;
	end
assign N11846 = x_reg_22__retimed_I7002_QOUT;
reg x_reg_22__retimed_I6999_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6999_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716;
	end
assign N11838 = x_reg_22__retimed_I6999_QOUT;
reg x_reg_22__retimed_I6996_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6996_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418;
	end
assign N11830 = x_reg_22__retimed_I6996_QOUT;
reg x_reg_22__retimed_I6993_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6993_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749;
	end
assign N11822 = x_reg_22__retimed_I6993_QOUT;
reg x_reg_22__retimed_I6990_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6990_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452;
	end
assign N11814 = x_reg_22__retimed_I6990_QOUT;
reg x_reg_22__retimed_I6987_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6987_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781;
	end
assign N11806 = x_reg_22__retimed_I6987_QOUT;
reg x_reg_22__retimed_I6984_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6984_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492;
	end
assign N11798 = x_reg_22__retimed_I6984_QOUT;
reg x_reg_22__retimed_I6981_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6981_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985;
	end
assign N11788 = x_reg_22__retimed_I6981_QOUT;
reg x_reg_11__retimed_I6955_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I6955_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896;
	end
assign N11722 = x_reg_11__retimed_I6955_QOUT;
reg x_reg_12__retimed_I6953_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I6953_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546;
	end
assign N11717 = x_reg_12__retimed_I6953_QOUT;
reg x_reg_13__retimed_I6951_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I6951_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813;
	end
assign N11712 = x_reg_13__retimed_I6951_QOUT;
reg x_reg_14__retimed_I6949_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I6949_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465;
	end
assign N11707 = x_reg_14__retimed_I6949_QOUT;
reg x_reg_15__retimed_I6947_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I6947_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735;
	end
assign N11702 = x_reg_15__retimed_I6947_QOUT;
reg x_reg_16__retimed_I6945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I6945_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006;
	end
assign N11697 = x_reg_16__retimed_I6945_QOUT;
reg x_reg_17__retimed_I6943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I6943_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654;
	end
assign N11692 = x_reg_17__retimed_I6943_QOUT;
reg x_reg_18__retimed_I6941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I6941_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929;
	end
assign N11687 = x_reg_18__retimed_I6941_QOUT;
reg x_reg_19__retimed_I6939_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I6939_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580;
	end
assign N11682 = x_reg_19__retimed_I6939_QOUT;
reg x_reg_20__retimed_I6937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I6937_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983;
	end
assign N11677 = x_reg_20__retimed_I6937_QOUT;
reg x_reg_21__retimed_I6935_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I6935_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503;
	end
assign N11672 = x_reg_21__retimed_I6935_QOUT;
reg x_reg_22__retimed_I6933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6933_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772;
	end
assign N11667 = x_reg_22__retimed_I6933_QOUT;
reg x_reg_22__retimed_I6864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6864_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29;
	end
assign N11506 = x_reg_22__retimed_I6864_QOUT;
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7517 (.Y(N13149), .A(N11506));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7518 (.Y(N13150), .A(N13149));
reg x_reg_22__retimed_I6863_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6863_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67;
	end
assign N11504 = x_reg_22__retimed_I6863_QOUT;
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7573 (.Y(N13151), .A(N11504));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7524 (.Y(N13156), .A(N13151));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7523 (.Y(N13155), .A(N13151));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7522 (.Y(N13154), .A(N13151));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7521 (.Y(N13153), .A(N13151));
reg x_reg_22__retimed_I6861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I6861_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
	end
assign N11500 = x_reg_22__retimed_I6861_QOUT;
INVX3 float_div_cynw_cm_float_rcp_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353), .A(a_exp[7]), .B(a_exp[0]));
AND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I2 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL float_div_cynw_cm_float_rcp_E8_M23_4_I3 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743), .A(a_exp[6]), .B(a_exp[5]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I4 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I5 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I6 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I8 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I9 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I10 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I11 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I12 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .A(a_man[18]), .B(a_man[17]));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I13 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I14 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B(a_man[16]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408), .D(a_man[15]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I15 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I16 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I17 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I18 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I19 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I20 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I21 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_rcp_E8_M23_4_I22 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I23 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I24 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .A(a_exp[1]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I25 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]), .A(a_exp[0]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I26 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I27 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I28 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I29 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .A(a_exp[3]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I30 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457), .A(a_exp[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I31 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I32 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .A(a_exp[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I33 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I34 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I35 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_4_I36 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I37 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I38 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I39 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .A(a_exp[7]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I40 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444), .A(a_exp[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I41 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I42 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I43 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .A(a_exp[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I44 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464));
NOR4BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I45 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I46 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I47 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8]));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I48 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I49 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
OR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I50 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I51 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I52 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I53 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A(a_man[22]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I54 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A(a_man[21]));
CLKINVX6 float_div_cynw_cm_float_rcp_E8_M23_4_I55 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I56 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I57 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .B(a_man[20]));
INVX3 float_div_cynw_cm_float_rcp_E8_M23_4_I58 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A(a_man[20]));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_4_I59 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A(a_man[18]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I60 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .A(a_man[16]), .B(a_man[17]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I61 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I62 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I63 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I64 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071), .B1(a_man[21]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I65 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .A(a_man[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I66 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .A(a_man[16]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I67 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I68 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I69 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I70 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I71 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I72 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I73 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I74 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I75 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I76 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .A(a_man[17]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I77 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I78 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I79 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I80 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I81 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I82 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .A(a_man[17]), .B(a_man[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I83 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I84 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .A1N(a_man[19]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I85 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I86 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I87 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I88 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I89 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I90 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I91 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I92 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I93 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I94 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I95 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I96 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I97 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I98 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I99 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809), .B1(a_man[21]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022), .B0(a_man[19]), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054), .A(a_man[19]), .B(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415), .B1(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I109 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841), .A(1'B0), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I110 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213), .B1(a_man[22]));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .A(a_man[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .A0(a_man[16]), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I151 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I155 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I161 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I162 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I163 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I164 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I165 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945), .B1(a_man[22]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783), .A(1'B1), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I167 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I169 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I170 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I171 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .A(a_man[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I173 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400), .B1(a_man[20]));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I199 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I201 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589), .A1N(a_man[21]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .A(a_man[14]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .A(a_man[13]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I207 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I211 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I213 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I214 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I215 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I217 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I221 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603), .B0(a_man[18]), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I223 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I225 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I227 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637), .A(a_man[12]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_4_I242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848), .B(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I253 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888), .A(a_man[11]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_4_I256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I259 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I269 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I271 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I272 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I273 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I274 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I275 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I276 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .A(a_man[10]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I302 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I303 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I304 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I305 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I310 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I314 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I318 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I319 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I323 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I324 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I325 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I326 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I327 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I328 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I329 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I348 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I349 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I350 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I351 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747), .A(a_man[9]));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_4_I355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I371 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I372 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I373 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I377 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I378 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648), .A(a_man[8]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I384 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I387 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I388 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I389 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I390 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I391 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I392 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I393 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .A(a_man[7]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I423 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I424 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I428 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I432 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I433 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I439 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I440 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I444 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I445 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I446 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I448 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I449 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I450 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B0(a_man[18]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I471 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I472 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I473 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I474 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I475 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I476 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .A(a_man[6]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I481 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I485 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I486 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430), .A(a_man[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I490 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I495 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I496 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I497 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I498 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I499 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I500 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I501 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I502 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I503 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I504 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I505 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I506 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I507 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I520 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I525 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B(a_man[18]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I526 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I541 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I542 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I543 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I547 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698), .A(a_man[5]));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I548 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698));
INVX2 float_div_cynw_cm_float_rcp_E8_M23_4_I549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I552 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I571 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I573 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I575 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I576 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I577 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I578 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I579 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I580 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I581 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I582 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I584 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I585 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I587 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I588 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I589 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I592 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I594 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I598 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I606 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I608 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I612 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I613 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I614 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I616 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I618 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .A(a_man[4]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .A(a_man[3]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I640 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I641 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I645 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I646 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I650 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I654 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I666 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I671 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I672 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I677 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I679 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I681 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I682 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I686 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I690 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I691 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I692 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I693 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I694 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I695 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I696 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I697 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I698 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I706 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I707 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I708 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I710 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I711 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I712 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I713 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I714 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I715 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I719 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I723 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I724 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I725 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I726 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I729 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I730 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I733 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .A(a_man[2]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I734 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .A(a_man[0]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .A(a_man[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I736 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I737 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I738 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I741 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I742 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I746 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I747 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I748 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I749 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I750 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I751 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I752 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I753 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I757 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .A(a_man[22]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I759 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I760 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I763 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2801), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2821), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2600));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I767 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I768 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I769 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7737 (.Y(N13667), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7738 (.Y(N13630), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7739 (.CO(N13649), .S(N13639), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7740 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663), .S(N13661), .A(N13667), .B(N13630), .CI(N13649));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I783 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I786 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I789 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I790 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I795 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I796 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I798 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I799 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I800 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I801 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I802 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I803 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2686), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2581), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2717));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I807 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I808 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I809 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I810 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2617));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I811 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I812 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I813 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I814 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I816 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I817 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I818 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I819 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I825 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7711 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614), .S(N13556), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I827 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I833 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I834 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I835 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I836 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I839 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I841 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7712 (.CO(N13590), .S(N13579), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7713 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754), .S(N13550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587), .CI(N13590));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I844 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I845 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I846 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I850 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I851 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I852 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I855 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7714 (.CO(N13583), .S(N13570), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2677), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7715 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .S(N13542), .A(N13583), .B(N13556), .CI(N13550));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I860 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I861 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I862 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I868 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I869 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I870 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I871 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7680 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702), .S(N13440), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I873 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7681 (.CO(N13474), .S(N13459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7682 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846), .S(N13486), .A(N13474), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I881 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I886 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I887 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7683 (.CO(N13466), .S(N13452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7684 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .S(N13478), .A(N13440), .B(N13466), .CI(N13486));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I890 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I891 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I892 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I893 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I894 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I898 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I899 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I900 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I905 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I913 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I914 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7692 (.CO(N13445), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I918 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I919 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I920 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I921 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I922 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I923 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I924 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I925 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I926 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7685 (.CO(N13457), .S(N13447), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7686 (.CO(N13484), .S(N13472), .A(N13457), .B(N13459), .CI(N13452));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7687 (.Y(N13443), .A(N13484));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7688 (.Y(N13468), .A(N13443));
MXI2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7689 (.Y(N13479), .A(N13468), .B(N13443), .S0(N13478));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7690 (.CO(N13464), .S(N13450), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726), .CI(N13447));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7691 (.Y(N13476), .A(N13464), .B(N13472));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7693 (.Y(N13455), .A(N13445), .B(N13450));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7694 (.Y(N13470), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797));
OAI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7695 (.Y(N13482), .A0(N13445), .A1(N13450), .B0(N13455), .B1(N13470));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7696 (.Y(N13461), .A(N13472));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7697 (.Y(N13436), .A(N13464));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7698 (.Y(N13463), .A0(N13461), .A1(N13436), .B0(N13476), .B1(N13482));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7699 (.Y(N13460), .A(N13484), .B(N13478));
OAI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576), .A0(N13463), .A1(N13479), .B0(N13460));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I933 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7716 (.CO(N13577), .S(N13564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7717 (.CO(N13548), .S(N13588), .A(N13579), .B(N13577), .CI(N13570));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795), .A(N13548), .B(N13542));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7719 (.CO(N13581), .S(N13568), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2608), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2760), .CI(N13564));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652), .A(N13581), .B(N13588));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7721 (.Y(N13553), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583), .B(N13568));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7722 (.Y(N13562), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11756), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11758));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7723 (.Y(N13575), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2583), .B(N13568));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7724 (.Y(N13557), .A0(N13553), .A1(N13562), .B0(N13575));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7725 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871), .A0(N13553), .A1(N13562), .B0(N13575));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7726 (.Y(N13571), .A(N13588));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7727 (.Y(N13543), .A(N13581));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7728 (.Y(N13546), .A(N13581), .B(N13588));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7729 (.Y(N13586), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652), .B(N13557));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7730 (.Y(N13573), .A(N13546), .B(N13586));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749), .A0(N13571), .A1(N13543), .B0(N13586));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7732 (.Y(N13566), .A(N13548), .B(N13542));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7733 (.Y(N13551), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795), .B(N13573));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7734 (.Y(N13591), .A(N13566), .B(N13551));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7735 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .A(N13591));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I943 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2758));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2828));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I947 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2835), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2858));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7741 (.CO(N13642), .S(N13634), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7742 (.Y(N13655), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7743 (.CO(N13628), .S(N13665), .A(N13642), .B(N13655), .CI(N13639));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813), .A(N13661), .B(N13628));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7745 (.CO(N13659), .S(N13647), .A(N13634), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2649), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2792));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7746 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667), .A(N13659), .B(N13665));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852), .A(N13647), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2641));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7749 (.Y(N13653), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2606), .B(N13647));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7750 (.Y(N13636), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .B0(N13653));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7751 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .B0(N13653));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7752 (.Y(N13650), .A(N13665));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7753 (.Y(N13671), .A(N13659));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7754 (.Y(N13626), .A(N13665), .B(N13659));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7755 (.Y(N13663), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667), .B(N13636));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7756 (.Y(N13651), .A(N13626), .B(N13663));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7757 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601), .A0(N13650), .A1(N13671), .B0(N13663));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7758 (.Y(N13645), .A(N13661), .B(N13628));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7759 (.Y(N13632), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813), .B(N13651));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7760 (.Y(N13668), .A(N13645), .B(N13632));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634), .A(N13668));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I955 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2734), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2663));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7704 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7705 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2881));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7706 (.Y(N13530), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I7707 (.Y(N13518), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811), .B0(N13530));
NAND2BXL float_div_cynw_cm_float_rcp_E8_M23_4_I7708 (.Y(N13521), .AN(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7709 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176), .A(N13521), .B(N13518));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I963 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I964 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I965 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I966 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I967 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I968 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I974 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I975 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I979 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I983 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I984 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I985 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I986 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I987 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798), .B(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I992 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
CLKXOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I993 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769));
BUFX2 float_div_cynw_cm_float_rcp_E8_M23_4_I994 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I995 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I996 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I997 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1001 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1003 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1004 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1005 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917), .A(a_man[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1006 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1009 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010), .A(N12087), .B(N12085), .CI(N12089));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1012 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .A(a_man[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1013 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1014 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1018 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1019 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1020 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1021 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1023 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1024 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1025 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1026 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1030 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1033 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1034 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1035 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1036 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1040 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1043 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1045 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1046 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1047 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1048 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1049 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1050 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1051 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1054 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1055 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1057 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1058 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1059 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1060 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1061 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1062 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1063 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1067 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1068 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1069 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1070 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1071 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1072 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1073 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1077 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1078 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1079 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1080 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .A(a_man[16]), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1081 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1085 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1087 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1088 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1089 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1090 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1095 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1096 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1097 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1098 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1099 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1104 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1105 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1108 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1110 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1111 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1113 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1114 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1117 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1118 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1120 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1122 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542), .B1(a_man[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1125 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1136 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1140 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1145 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1146 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1147 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1151 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1152 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1153 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1154 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1155 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1156 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1157 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1159 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1160 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1161 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1162 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1163 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1164 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1165 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1166 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1167 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1168 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1169 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1170 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1172 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7630 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722), .S(N13370), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530), .B(N12003), .CI(N12007));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1173 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722), .B(N11937), .CI(N11941));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1175 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1183 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064), .B1(a_man[21]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1185 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1187 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1189 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1190 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1192 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1193 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1198 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1199 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1200 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1201 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1202 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1203 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1205 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1207 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1209 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1211 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1213 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1215 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1216 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1217 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1219 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1220 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1221 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1222 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1223 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1224 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1225 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1226 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7631 (.CO(N13400), .S(N13391), .A(N12042), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010), .CI(N12044));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7632 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589), .S(N13364), .A(N13400), .B(N11966), .CI(N13370));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1229 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1231 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1233 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1235 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1237 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1239 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1241 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1243 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1254 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1255 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1256 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1257 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1258 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1259 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1260 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1261 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1262 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1263 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1264 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1265 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1266 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105), .B1(a_man[21]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1267 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1268 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1269 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1270 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1271 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1272 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]), .A(N12240), .B(N12238), .CI(N12242));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1274 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1275 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1276 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1277 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1278 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1279 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1281 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1282 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1283 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1284 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1285 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1286 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1287 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1288 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1289 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1290 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1291 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1292 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1293 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1294 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1295 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1296 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1297 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1298 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1299 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1300 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1301 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1302 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1303 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1304 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1305 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1306 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1307 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1308 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1309 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1310 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1311 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1312 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1313 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1314 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1315 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1316 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1317 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1318 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1319 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1320 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1321 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1322 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1323 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1324 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1325 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1326 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1327 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1328 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1329 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1330 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1331 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1332 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1333 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1334 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1335 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1336 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1337 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1338 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1339 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1340 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1341 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1342 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1343 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1344 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1345 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1346 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1347 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1348 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552), .A(N12177), .B(N12175), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1352 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1353 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1354 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1355 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1356 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1357 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1358 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1359 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1360 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737), .B1(a_man[20]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1361 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904), .A(a_man[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1362 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1363 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1364 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1365 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1366 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1367 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1368 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1369 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1370 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1371 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1372 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1373 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1374 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1375 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1376 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1377 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111), .B1(a_man[20]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1378 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1379 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1380 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1381 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1382 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1383 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1384 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1385 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1386 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1387 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1388 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1389 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1390 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1391 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1392 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]), .A(N12295), .B(N12293), .CI(N12297));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1393 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817), .A(N12183), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1394 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1395 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985), .B1(a_man[19]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1396 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1397 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1398 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1399 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1400 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1401 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1402 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1403 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1404 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1405 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1406 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1407 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1408 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1409 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B0(a_man[17]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1410 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1411 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1412 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1413 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264), .B1(a_man[22]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1414 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1415 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1416 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1417 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1418 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1419 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1420 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1421 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1422 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1423 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1424 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1425 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1426 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1427 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1428 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1429 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1430 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1431 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1432 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1433 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1434 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1435 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1436 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1437 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1438 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1439 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1440 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1441 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1442 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1443 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1444 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1445 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1446 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1447 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1448 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1449 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1450 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(a_man[16]), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1451 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1452 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1453 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1454 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1455 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1456 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1457 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1458 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1459 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1460 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1461 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1462 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1463 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1464 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1465 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1466 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1467 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1468 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1469 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1470 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1471 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1472 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817), .B(N12122), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1475 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1476 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1477 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1478 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1479 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1480 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1481 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1482 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1483 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1484 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1485 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1486 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1487 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1488 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1489 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1490 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1491 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1492 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1493 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1494 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1495 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1496 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1497 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1498 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1499 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1500 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1501 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1502 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1503 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1504 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1505 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1506 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[18]), .B0(a_man[16]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1507 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1508 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1509 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1510 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1511 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1512 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1513 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1514 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B1(a_man[19]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1515 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(a_man[17]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1516 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1517 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1518 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1519 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1520 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1521 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1522 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1523 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1524 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1525 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1526 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1527 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1528 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1529 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1530 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1531 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1532 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1533 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1534 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1535 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1536 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1537 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1538 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1539 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1540 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1541 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1542 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1543 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1544 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1545 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1546 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1547 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1548 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1549 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1550 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1551 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1552 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1553 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1554 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1555 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1556 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1557 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1558 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1559 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1560 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1561 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1562 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1564 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1565 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1566 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1567 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1568 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1569 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1570 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1571 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1572 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1573 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1574 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1575 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1576 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1578 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1579 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1580 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1581 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299), .A(N12445), .B(N12443), .CI(N12447));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1582 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1583 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376), .B(N12285), .CI(N12289));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1584 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1585 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868), .A(N12169), .B(N12167), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1586 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1588 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1589 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1590 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1591 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1592 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1593 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1594 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1596 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1597 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1598 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1599 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1600 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1601 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1602 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1605 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1606 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1607 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1608 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1609 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1610 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1611 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1612 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1613 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1614 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1615 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1616 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1617 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1619 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1620 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1621 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1623 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1624 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1626 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1627 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1629 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1630 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1631 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1632 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1633 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1634 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1635 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1636 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1637 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1638 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1639 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1640 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1641 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1645 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1646 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1648 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1649 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1650 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1652 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1653 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1654 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1655 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1656 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1657 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1658 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1659 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1660 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1661 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1662 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1663 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1664 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1665 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1666 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1667 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1668 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1669 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1670 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1671 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1672 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1673 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1674 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1675 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1676 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1677 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1678 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1679 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1680 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1681 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1682 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1683 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1684 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1685 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1686 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1687 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889), .B1(a_man[20]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1688 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1689 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1690 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1691 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1692 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218), .B1(a_man[22]));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I1693 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1694 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1695 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1696 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1697 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1698 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1699 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1700 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1701 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1702 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1703 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1704 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1705 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1706 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1707 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370), .A(N12506), .B(N12504), .CI(N12508));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1708 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1709 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239), .A(N12512), .B(N12516), .CI(N12514));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1710 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104), .B(N12435), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1711 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312), .B(N12383), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1712 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7588 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557), .S(N13256), .A(N12220), .B(N12218), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7589 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497), .S(N13281), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1715 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1716 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1717 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1718 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1719 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1720 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1721 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1722 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1723 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1724 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1725 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1726 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1727 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1728 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1729 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1730 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1731 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1732 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1733 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1734 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1735 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1736 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1737 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1738 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1739 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1740 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1741 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1742 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1743 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1744 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1745 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1746 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1747 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1748 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1749 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1750 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1751 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1752 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1753 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1754 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1755 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1756 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1757 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7590 (.CO(N13259), .S(N13248), .A(N12279), .B(N12277), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7591 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .S(N13273), .A(N13259), .B(N13281), .CI(N13256));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1760 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1761 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1762 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1763 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1764 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1765 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1766 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1767 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1768 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1769 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1770 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1771 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1772 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1773 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1774 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1775 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1776 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1777 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1778 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1779 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1780 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1781 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1782 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1783 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1784 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1785 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1786 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1787 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1788 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1789 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1790 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1791 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1792 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1793 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1794 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1795 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1796 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1797 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1798 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1799 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1800 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1801 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1802 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1803 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1804 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1805 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1806 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1807 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1808 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1809 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1810 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1811 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1812 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1813 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1814 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1815 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]), .A(N12423), .B(N12421), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1820 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1821 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1822 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1823 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1824 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1825 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1826 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1827 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1828 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1829 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1830 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1831 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1832 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1833 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1834 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1835 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1836 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1837 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009), .B1(a_man[22]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1838 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1839 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1840 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1841 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1842 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1843 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1844 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1845 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1846 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1847 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1848 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1849 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1850 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1851 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1852 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1853 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1854 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1855 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1856 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1857 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1858 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1859 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1860 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1861 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1862 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1863 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1864 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1865 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1866 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1867 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1868 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1869 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1870 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1871 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1872 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1873 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1874 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1875 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1876 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1877 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1878 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1879 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1880 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1881 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1882 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1883 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1884 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1885 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1886 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1887 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1888 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1889 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1890 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1891 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1892 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_4_I1893 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1894 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]), .A(N12490), .B(N12488), .CI(N12492));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1895 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675), .A(N12429), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1896 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655), .A(N12365), .B(N12363), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1897 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]), .A(N12498), .B(N12496), .CI(N12500));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1898 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I1901 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1902 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[17]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1903 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1904 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1905 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1906 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1907 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1908 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1909 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1910 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1911 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1912 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1913 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641), .A1(a_man[16]), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036), .B1(a_man[18]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1914 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1915 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600), .B1(a_man[19]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1916 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836), .B1(a_man[20]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1917 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474), .B1(a_man[21]));
AOI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I1918 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812), .B1(a_man[22]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1919 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1920 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1921 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1922 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1923 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1924 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763), .A(N12415), .B(N12413), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1925 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1927 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1928 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1929 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1930 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1931 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1932 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1933 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1934 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1935 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1936 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1937 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]), .A(N12552), .B(N12550), .CI(N12554));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1938 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861), .A(N12482), .B(N12480), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1939 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1940 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1941 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1942 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1943 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1944 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1945 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1946 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1947 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1948 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1949 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1950 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1951 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1952 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1953 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1954 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1955 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1956 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1957 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1958 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1959 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1960 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1961 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1962 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1963 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1964 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1965 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1966 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1967 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964), .A(N12544), .B(N12542), .CI(N12627));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1968 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1969 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1970 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1971 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1972 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1973 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1974 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1975 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1976 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1977 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1978 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1979 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1980 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1981 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1982 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1983 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1984 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1985 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1986 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1987 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1988 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1989 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1990 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1991 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1992 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1993 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1994 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1995 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1996 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442), .A(N12580), .B(N12578), .CI(N12582));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I1997 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1998 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I1999 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2000 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2001 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2002 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2003 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2004 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2005 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2006 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2007 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2008 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2009 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2010 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2011 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2012 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2013 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2014 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545), .A(N12529), .B(N12625), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2015 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2016 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2017 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2018 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2019 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2020 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2021 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2022 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2023 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2024 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2025 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2026 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2027 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2028 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2029 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2030 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2031 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2032 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2033 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2034 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2035 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2036 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2037 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2038 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2039 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2040 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2041 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2042 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2043 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2044 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2045 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2046 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2047 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2048 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2049 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2050 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971), .A(N12607), .B(N12605), .CI(N12609));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2051 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761), .A(N12562), .B(N12560), .CI(N12564));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2052 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2053 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2054 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2055 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2056 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2057 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2058 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2059 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2060 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2061 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2062 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2063 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2064 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2065 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2066 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2067 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2068 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2069 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2070 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2071 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2072 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2073 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826), .A(N12567), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2074 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2075 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2076 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2077 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2078 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2079 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2080 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2081 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2082 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2083 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2084 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2085 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2086 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2087 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2088 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2089 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2090 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2091 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2092 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2093 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2094 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2095 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2096 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2097 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2098 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2099 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2100 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2101 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2102 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2103 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2104 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2105 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2106 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2107 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2108 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2109 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2110 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2111 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2112 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2113 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2114 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2115 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2116 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2117 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2118 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2119 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2120 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2121 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2122 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]));
AND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2123 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2124 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2125 (.CO(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .S(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2126 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823));
NOR4X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2127 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533), .D(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2128 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2129 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2130 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2131 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2132 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2133 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2134 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2135 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2136 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2137 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2138 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2139 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2140 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948), .A0(N12591), .A1(N12585), .B0(N12587), .B1(N12589));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2141 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699), .A(N12567), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971));
AOI21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2142 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699));
OAI22XL float_div_cynw_cm_float_rcp_E8_M23_4_I2143 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2144 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2145 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545));
AO21XL float_div_cynw_cm_float_rcp_E8_M23_4_I2146 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615));
AOI2BB2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7279 (.Y(N12613), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7280 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558), .A(N12613));
OAI2BB2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2148 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733));
OAI2BB2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2149 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869), .B1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2150 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927));
ADDHX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7592 (.CO(N13254), .S(N13241), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7593 (.CO(N13279), .S(N13263), .A(N12327), .B(N12325), .CI(N13241));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7594 (.CO(N13246), .S(N13236), .A(N13254), .B(N13279), .CI(N13248));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7595 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593), .A(N13246), .B(N13273));
ADDFXL float_div_cynw_cm_float_rcp_E8_M23_4_I7596 (.CO(N13229), .S(N13271), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578), .CI(N13263));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7597 (.Y(N13274), .A(N13229));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7598 (.Y(N13251), .A(N13274), .B(N13236));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7599 (.Y(N13232), .A(N13251));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7600 (.Y(N13266), .A(N13229));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7601 (.Y(N13238), .A(N13266), .B(N13236));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7602 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940), .A(N13236), .B(N13229));
CLKXOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7603 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .B(N13271));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7604 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7605 (.Y(N13277), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439), .B(N13271));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7606 (.Y(N13234), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7607 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668), .B0(N13277));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7608 (.Y(N13242), .A(N13236));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7609 (.Y(N13264), .A(N13229), .B(N13236));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7610 (.Y(N13269), .A0(N13238), .A1(N13232), .B0(N13277), .B1(N13234));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7611 (.Y(N13250), .A(N13269));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7612 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500), .A0N(N13242), .A1N(N13274), .B0(N13250));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7613 (.Y(N13268), .A(N13246), .B(N13273));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7614 (.Y(N13267), .A0(N13264), .A1(N13269), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7615 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .A(N13268), .B(N13267));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2158 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2159 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2160 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7633 (.CO(N13395), .S(N13385), .A(N12132), .B(N12130), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7634 (.CO(N13368), .S(N13353), .A(N13385), .B(N12077), .CI(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7635 (.CO(N13389), .S(N13380), .A(N13368), .B(N13395), .CI(N13391));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7636 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704), .A(N13364), .B(N13389));
ADDFX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7637 (.CO(N13373), .S(N13362), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957), .CI(N13353));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7638 (.Y(N13371), .A(N13380));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7639 (.Y(N13376), .A(N13373), .B(N13371));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7640 (.Y(N13356), .A(N13373));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7641 (.Y(N13382), .A(N13380), .B(N13356));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7642 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430), .A(N13373), .B(N13380));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7643 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782), .A(N13362), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7644 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7645 (.Y(N13366), .A(N13362), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7646 (.Y(N13378), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7647 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .B0(N13366));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7648 (.Y(N13354), .A(N13373), .B(N13380));
AOI22X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7649 (.Y(N13360), .A0(N13382), .A1(N13376), .B0(N13366), .B1(N13378));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7650 (.Y(N13392), .A(N13360));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7651 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996), .A0N(N13371), .A1N(N13356), .B0(N13392));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7652 (.Y(N13359), .A(N13364), .B(N13389));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7653 (.Y(N13358), .A0(N13354), .A1(N13360), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7654 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .A(N13359), .B(N13358));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2168 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2172 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2174 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568));
XOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7617 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623), .A(N11886), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7618 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .B0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7619 (.Y(N13337), .A(N11886), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7620 (.Y(N13329), .A(N13337));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7621 (.Y(N13319), .A0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .B0(N13329));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7622 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .A0N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .B0(N13337));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7623 (.Y(N13318), .A(N11722));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7624 (.Y(N13326), .A(N13318), .B(N13319));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7625 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567), .A0N(N11722), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .B0(N11862));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7626 (.Y(N13322), .A(N11862));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7627 (.Y(N13330), .A0(N13322), .A1(N13326), .B0(N11717));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7628 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .A(N11854), .B(N13330));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2176 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2177 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .A0N(N11712), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .B0(N11846));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2178 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2179 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .A0N(N11707), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .B0(N11838));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2180 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2181 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736), .A0N(N11702), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .B0(N11830));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2182 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2184 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2186 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2188 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7577 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .A0N(N11697), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736), .B0(N11822));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7578 (.Y(N13204), .A(N11814));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7579 (.Y(N13205), .A0(N11692), .A1(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .B0(N13204));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7580 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588), .A0N(N11692), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .B0(N11814));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7581 (.Y(N13209), .A(N11687));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7582 (.Y(N13212), .A(N13209), .B(N13205));
OAI2BB1X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7583 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608), .A0N(N11687), .A1N(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588), .B0(N11806));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7584 (.Y(N13202), .A(N11806));
OAI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7585 (.Y(N13215), .A0(N13202), .A1(N13212), .B0(N11682));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7586 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899), .A(N11798), .B(N13215));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7281 (.Y(N12618), .AN(N11677), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2191 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7562 (.Y(N13167), .A(N11788));
INVX1 float_div_cynw_cm_float_rcp_E8_M23_4_I7563 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834), .A(N12618));
NAND2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7564 (.Y(N13180), .A(N11672), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7565 (.Y(N13172), .A(N11667));
AOI21X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7566 (.Y(N13181), .A0(N13167), .A1(N13180), .B0(N13172));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7567 (.Y(N13170), .A(N13167));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7568 (.Y(N13182), .A(N11672));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7569 (.Y(N13174), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834));
NOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7570 (.Y(N13166), .A(N13182), .B(N13174));
NOR3X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7571 (.Y(N13164), .A(N11667), .B(N13170), .C(N13166));
NAND2XL float_div_cynw_cm_float_rcp_E8_M23_4_I7572 (.Y(N13178), .A(N11500), .B(N11506));
OAI31X1 float_div_cynw_cm_float_rcp_E8_M23_4_I7574 (.Y(x[22]), .A0(N13164), .A1(N13181), .A2(N13151), .B0(N13178));
INVXL float_div_cynw_cm_float_rcp_E8_M23_4_I7575 (.Y(N13152), .A(N13151));
NOR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2194 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2195 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896), .B(a_man[22]));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2196 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2197 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2200 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834), .B(N11672));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2201 (.Y(x[21]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]), .S0(N13154));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2202 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899), .B(N11677));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2203 (.Y(x[20]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]), .S0(N13156));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2204 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608), .B(N11682));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2205 (.Y(x[19]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]), .S0(N13155));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2206 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588), .B(N11687));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2207 (.Y(x[18]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]), .S0(N13153));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2208 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831), .B(N11692));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2209 (.Y(x[17]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]), .S0(N13154));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2210 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736), .B(N11697));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2211 (.Y(x[16]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]), .S0(N13153));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2212 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911), .B(N11702));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2213 (.Y(x[15]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]), .S0(N13155));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2214 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728), .B(N11707));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2215 (.Y(x[14]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31]), .S0(N13155));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2216 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820), .B(N11712));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2217 (.Y(x[13]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]), .S0(N13154));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2218 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567), .B(N11717));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2219 (.Y(x[12]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]), .S0(N13152));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2220 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579), .B(N11722));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2221 (.Y(x[11]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]), .S0(N13152));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2222 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2223 (.Y(x[10]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]), .S0(N13152));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2224 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2225 (.Y(x[9]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]), .S0(N13154));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2226 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2227 (.Y(x[8]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]), .S0(N13156));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2228 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2229 (.Y(x[7]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]), .S0(N13155));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2230 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2231 (.Y(x[6]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]), .S0(N13153));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2232 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2233 (.Y(x[5]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]), .S0(N13153));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2234 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2235 (.Y(x[4]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]), .S0(N13153));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2236 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2237 (.Y(x[3]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]), .S0(N13155));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2238 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2239 (.Y(x[2]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]), .S0(N13156));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2240 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2241 (.Y(x[1]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]), .S0(N13154));
XNOR2X1 float_div_cynw_cm_float_rcp_E8_M23_4_I2242 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2243 (.Y(x[0]), .A(N13150), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]), .S0(N13152));
OR2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2244 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34));
NOR3XL float_div_cynw_cm_float_rcp_E8_M23_4_I2245 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34), .C(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2246 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2247 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2248 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2249 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2250 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2251 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2252 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
MX2XL float_div_cynw_cm_float_rcp_E8_M23_4_I2253 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23]), .A(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]), .S0(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42));
NOR2BX1 float_div_cynw_cm_float_rcp_E8_M23_4_I2254 (.Y(float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31]), .AN(a_sign), .B(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29));
reg x_reg_23__I2278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__I2278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23];
	end
assign x[23] = x_reg_23__I2278_QOUT;
reg x_reg_24__I2279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_24__I2279_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24];
	end
assign x[24] = x_reg_24__I2279_QOUT;
reg x_reg_25__I2280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_25__I2280_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25];
	end
assign x[25] = x_reg_25__I2280_QOUT;
reg x_reg_26__I2281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_26__I2281_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26];
	end
assign x[26] = x_reg_26__I2281_QOUT;
reg x_reg_27__I2282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_27__I2282_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27];
	end
assign x[27] = x_reg_27__I2282_QOUT;
reg x_reg_28__I2283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_28__I2283_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28];
	end
assign x[28] = x_reg_28__I2283_QOUT;
reg x_reg_29__I2284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__I2284_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29];
	end
assign x[29] = x_reg_29__I2284_QOUT;
reg x_reg_30__I2285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_30__I2285_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30];
	end
assign x[30] = x_reg_30__I2285_QOUT;
reg x_reg_31__I2286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I2286_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_31__I2286_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0] = x[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1] = x[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2] = x[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3] = x[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4] = x[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5] = x[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6] = x[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7] = x[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8] = x[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9] = x[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10] = x[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11] = x[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12] = x[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13] = x[13];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  s7n4TQ/fohs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



