/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:25:07 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_1 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979;
wire N6566,N6655,N6659,N6666,N6673,N6680,N6687 
	,N6694,N6701,N6708,N6715,N6722,N6725,N6732,N6739 
	,N6746,N6753,N6760,N6767,N6774,N6781,N6788,N6795 
	,N6802,N6814,N6819,N6835,N6842,N6845,N6850,N6855 
	,N6860,N6868,N6873,N6878,N6885,N6888,N6893,N6900 
	,N6903,N6908,N6910,N6913,N6918,N6920,N6923,N6925 
	,N6930,N6933,N6935,N6938,N6973,N6978,N6980,N6997 
	,N7000,N7004,N7006,N7024,N7029,N7031,N7034,N7039 
	,N7051,N7063,N7065,N7070,N7072,N7074,N7079,N7083 
	,N7088,N7090,N7095,N7097,N7099,N7104,N7136,N7138 
	,N7146,N7152,N7158,N7162,N7170,N7172,N7178,N7180 
	,N7184,N7192,N7194,N7199,N7201,N7203,N7209,N7217 
	,N7219,N7225,N7227,N7232,N7236,N7249,N7251,N7567 
	,N7575,N7642,N7646,N7652,N7924,N7925,N7926,N7927 
	,N7928,N8020;
EDFFHQX1 x_reg_9__retimed_I4910 (.Q(N7652), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4908 (.Q(N7646), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__retimed_I4907 (.Q(N7642), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_5__retimed_I4876 (.Q(N7575), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_14__retimed_I4873 (.Q(N7567), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4735 (.Q(N7251), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4734 (.Q(N7249), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4731 (.Q(N7236), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4729 (.Q(N7232), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4727 (.Q(N7227), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4726 (.Q(N7225), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4724 (.Q(N7219), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4723 (.Q(N7217), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4721 (.Q(N7209), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4720 (.Q(N7203), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4719 (.Q(N7201), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4718 (.Q(N7199), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4716 (.Q(N7194), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4715 (.Q(N7192), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4712 (.Q(N7184), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4711 (.Q(N7180), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4710 (.Q(N7178), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4708 (.Q(N7172), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4707 (.Q(N7170), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4704 (.Q(N7162), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4703 (.Q(N7158), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4701 (.Q(N7152), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4699 (.Q(N7146), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4696 (.Q(N7138), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4695 (.Q(N7136), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I4683 (.Q(N7104), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__retimed_I4681 (.Q(N7099), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__retimed_I4680 (.Q(N7097), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__retimed_I4679 (.Q(N7095), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__retimed_I4677 (.Q(N7090), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__retimed_I4676 (.Q(N7088), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I4674 (.Q(N7083), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I4672 (.Q(N7079), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I4670 (.Q(N7074), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I4669 (.Q(N7072), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I4668 (.Q(N7070), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__retimed_I4666 (.Q(N7065), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__retimed_I4665 (.Q(N7063), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_24__retimed_I4660 (.Q(N7051), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_10__retimed_I4655 (.Q(N7039), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_8__retimed_I4653 (.Q(N7034), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_12__retimed_I4652 (.Q(N7031), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_12__retimed_I4651 (.Q(N7029), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_14__retimed_I4649 (.Q(N7024), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__retimed_I4642 (.Q(N7006), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__retimed_I4641 (.Q(N7004), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__retimed_I4639 (.Q(N7000), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__retimed_I4638 (.Q(N6997), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I4631 (.Q(N6980), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I4630 (.Q(N6978), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I4628 (.Q(N6973), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_1__retimed_I4623 (.Q(N6938), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_3__retimed_I4622 (.Q(N6935), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_3__retimed_I4621 (.Q(N6933), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_2__retimed_I4620 (.Q(N6930), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_11__retimed_I4618 (.Q(N6925), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_11__retimed_I4617 (.Q(N6923), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I4616 (.Q(N6920), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I4615 (.Q(N6918), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_13__retimed_I4613 (.Q(N6913), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_15__retimed_I4612 (.Q(N6910), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_15__retimed_I4611 (.Q(N6908), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_10__retimed_I4609 (.Q(N6903), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_6__retimed_I4608 (.Q(N6900), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_8__retimed_I4605 (.Q(N6893), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_12__retimed_I4603 (.Q(N6888), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_5__retimed_I4602 (.Q(N6885), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_9__retimed_I4599 (.Q(N6878), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_4__retimed_I4597 (.Q(N6873), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_14__retimed_I4595 (.Q(N6868), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__retimed_I4592 (.Q(N6860), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__retimed_I4590 (.Q(N6855), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__retimed_I4588 (.Q(N6850), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I4586 (.Q(N6845), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_22__retimed_I4585 (.Q(N6842), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I4582 (.Q(N6835), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__retimed_I4578 (.Q(N6819), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_23__retimed_I4576 (.Q(N6814), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_21__retimed_I4571 (.Q(N6802), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_20__retimed_I4568 (.Q(N6795), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_17__retimed_I4565 (.Q(N6788), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_13__retimed_I4562 (.Q(N6781), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_12__retimed_I4559 (.Q(N6774), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_11__retimed_I4556 (.Q(N6767), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_10__retimed_I4553 (.Q(N6760), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_8__retimed_I4550 (.Q(N6753), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_6__retimed_I4547 (.Q(N6746), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_3__retimed_I4544 (.Q(N6739), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_2__retimed_I4541 (.Q(N6732), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_0__retimed_I4538 (.Q(N6725), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_19__retimed_I4537 (.Q(N6722), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_18__retimed_I4534 (.Q(N6715), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_16__retimed_I4531 (.Q(N6708), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_15__retimed_I4528 (.Q(N6701), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_14__retimed_I4525 (.Q(N6694), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_9__retimed_I4522 (.Q(N6687), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_7__retimed_I4519 (.Q(N6680), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_5__retimed_I4516 (.Q(N6673), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_4__retimed_I4513 (.Q(N6666), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_1__retimed_I4510 (.Q(N6659), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_1__retimed_I4508 (.Q(N6655), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63), .E(bdw_enable), .CK(aclk));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5043 (.Y(N7924), .A(N6655));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5044 (.Y(N7925), .A(N7924));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5045 (.Y(N7926), .A(N6655));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5046 (.Y(N7927), .A(N7926));
EDFFHQX1 x_reg_0__retimed_I4483 (.Q(N6566), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[0]), .E(bdw_enable), .CK(aclk));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I0 (.Y(bdw_enable), .A(astall));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643), .A(a_exp[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563), .A(b_exp[7]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682), .A(a_exp[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562), .A(b_exp[6]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561), .A(b_exp[5]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560), .A(b_exp[4]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650), .A(a_exp[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559), .A(b_exp[3]));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602), .A(a_exp[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558), .A(b_exp[2]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557), .A(b_exp[1]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614), .A(a_exp[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556), .A(b_exp[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594), .A(a_exp[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640), .A(a_exp[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687), .A(a_exp[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625), .A(a_exp[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674), .A(a_exp[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609), .A(a_exp[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659), .A(a_exp[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4627), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4603));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17569), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17576));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I46 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I47 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631));
AO21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I48 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17597), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17588));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I49 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I50 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I51 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864), .A(a_man[20]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I52 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931), .A(a_man[21]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4865), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I56 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4891));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I57 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796), .A(a_man[19]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I58 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I59 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884), .A(a_man[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I60 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I61 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4819));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I62 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817), .A(a_man[17]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901), .A(a_man[16]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I66 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4924));
NAND3BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I67 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4873));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I68 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922), .A(a_man[14]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I69 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I70 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839), .A(a_man[15]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I71 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I72 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4878), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I73 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791), .A(a_man[12]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854), .A(a_man[13]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4832), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4853));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829), .A(a_man[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893), .A(a_man[9]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4889), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807), .A(a_man[10]));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875), .A(a_man[11]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875));
AOI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919), .A0N(b_man[10]), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4836), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4824));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847), .A(a_man[6]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912), .A(a_man[7]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4841), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934), .A(a_man[5]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866), .A(a_man[4]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4794));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4814));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338), .A(a_man[2]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801), .A(a_man[3]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4898), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911), .A(b_man[0]));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820), .A(a_man[1]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820));
OAI31X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914), .A0(a_man[0]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4800), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4835));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4933), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4846), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4880));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4881), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4914), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4848));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4828), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4927));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4790), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4874), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4823));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4899), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4935), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4868));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4923), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4856));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4921), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4837), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4869));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4882), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4816), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4915));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4802), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4919), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4888));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4929), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4863), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4810));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4825), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4910), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4857));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4789), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4822), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4906));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4908), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4792), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4876));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4938), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4818), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4903));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4871), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4805), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4904));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4917), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4851), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4799));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4806), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4926));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4897), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4812), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4845));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4861), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4859), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4830));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4928), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4809), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4894));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17571), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17578), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17586));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17595));
NAND2X8 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17590), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17580));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I156 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6017));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I157 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I158 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I159 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I160 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4671), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4656), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4619));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I161 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I162 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I163 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4645));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4595));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17592), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17583));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I166 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N567), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I167 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I168 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4677));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I172 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4630));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N566), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I176 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4614));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4666), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4594), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4640));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4658), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I180 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I181 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4592), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4667));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17869), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17859), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4647), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4680), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4621));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4611), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4685), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4626));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N569), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4602));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4650), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4687), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4625));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4688), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4668));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4684), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4682));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4649), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4634), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4638), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4607));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4623));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5094), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N572), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4654));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4641), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4631), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4615));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4637), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4609), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4635));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4601), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4695), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4610), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4673));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4613), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4661));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N571), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4606));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4596), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4692), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4678));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4598), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4697));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4648), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4662), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4624));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4591));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N570), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[5]));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5114), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5119), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5123));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17818), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17825));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17830), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17805));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17391));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233), .A(b_man[14]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5233), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206), .A(b_man[13]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5206), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4617), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4690));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556));
MXI2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N565), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[8]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249), .A(b_man[10]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5249), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222), .A(b_man[9]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5222), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
CLKINVX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[2]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164), .A(b_man[16]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5164), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259), .A(b_man[15]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5259), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180), .A(b_man[12]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5180), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153), .A(b_man[11]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5153), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
BUFX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[1]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141), .A(b_man[6]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5141), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237), .A(b_man[5]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5237), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433), .A(b_man[2]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253), .A(b_man[1]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5253), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195), .A(b_man[8]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5195), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168), .A(b_man[7]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5168), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210), .A(b_man[4]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5210), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184), .A(b_man[3]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5184), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[3]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201), .A(b_man[22]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5201), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4843), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175), .A(b_man[21]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5175), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217), .A(b_man[18]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5217), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191), .A(b_man[17]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148), .A(b_man[20]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5148), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244), .A(b_man[19]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5244), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480));
BUFX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[4]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[27]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[27]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N656), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[2]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655), .A(a_man[0]), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224), .A(a_man[0]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4911), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[26]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10782));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5355), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5387), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5548), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5420), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5363), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5541), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5574), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5482), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17372));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17371), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5551), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5583), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5492), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5366));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5558), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5454));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5519), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5486), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17895));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5431), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[24]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5555));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5429), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5490), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[2]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5529));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5495), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5527), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5471), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5397));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5559));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
NOR2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[5]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[2]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[5]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[8]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5415));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5447));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5569), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5383), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[16]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5922), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5901));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5899));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[10]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5521));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5581), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5441), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5503), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5401), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5474), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5434), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5464), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5375), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[23]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5568));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5518), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5577), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5359), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5563), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5480), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5545), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[19]));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5931), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5919));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17814), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17808));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5443), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5473), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5418), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5505));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
NOR2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[4]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445));
NOR2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[3]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5390));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5525), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5385), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5428), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5395), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5346));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5367), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5412), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5560));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5571), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[22]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[9]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5467));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5424));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5352), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5461), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5416), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5377), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[12]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5531));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5409), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5515), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5468), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5485), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5336));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5459), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5523), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5345), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[14]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5926), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5892));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5894), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5890));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[0]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5562));
NOR2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[6]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5554));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5499));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[1]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[1]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5506), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5406), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5498), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5538), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5398), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5496));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5350), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5445), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[20]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5905), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5909));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[7]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5357));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5391));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5513), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5578), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17945), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5452), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5373), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5438), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5423), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10862), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405));
OR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[15]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[17]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5916), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5924));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17821), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17828));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17835), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17811), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17829));
NAND3BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[1]));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6374), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5536), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5382), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[28]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[28]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N657));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6295));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6262), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5340), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5436), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[29]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[29]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6222));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I495 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6387));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[4]));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6477), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5396), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5489), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[30]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17952));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N659), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[5]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6364));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6254), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6179), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6394), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6325));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6336), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6474));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6211));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6365), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6467), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6293), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6201), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5450));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I527 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[31]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5544), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[31]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[31]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[31]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N660), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[6]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6249));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6355));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I535 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6177));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6281), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6435), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6475), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5504), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[32]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5348), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[32]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17959));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[7]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312));
XOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6462));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I549 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I550 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[34]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5458));
XNOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I552 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[34]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I553 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[9]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5365));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[33]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5405), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[33]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[33]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[33]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6465));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I564 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6176), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6459));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I566 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[8]));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6392), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6432), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6235), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I572 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6167), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6323), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6424), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6312), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6240));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6252), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6291), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I578 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I579 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6349));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I582 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I583 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6273));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I584 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6367), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6437));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I585 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6158));
INVXL buf1_A_I5091 (.Y(N8020), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17393));
INVXL buf1_A_I5092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955), .A(N8020));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__44));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I589 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I590 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I591 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[44]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5362));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[44]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[19]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[43]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5501));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[43]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I601 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5394));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[42]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I607 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[41]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5338));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I608 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[41]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I610 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[40]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5534));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I612 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[40]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I614 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[39]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5479), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[39]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I620 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I621 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[38]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[38]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I623 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I624 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I625 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[37]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5372));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I627 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[37]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I629 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I630 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[36]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5567));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I631 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[36]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I632 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I633 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[35]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5511));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[35]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I639 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I640 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I641 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6422));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6463));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I644 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[10]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I645 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6353), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I647 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6390), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I648 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I649 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[12]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I650 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[13]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[14]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[15]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17769), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17778));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[17]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[18]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I661 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6327), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6256));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6436), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6375), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6366));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6412), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6476));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I673 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6452));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6279));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6321));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6268), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6381), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6195));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6209), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I680 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6250), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6180), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6439));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6294), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6304), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6223));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I690 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6198), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6334));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I691 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I692 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I693 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5579));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I694 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[46]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I695 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I696 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[21]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I697 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I698 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I699 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5470));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I700 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[45]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I701 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6217));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6300));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I706 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6380));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6419));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6341), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6310), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6267));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6350), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6260), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6184));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[20]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I713 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I714 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6472), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I715 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I716 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6282), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6213));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6393), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6189), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6324));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6186), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6434));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6247));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6400));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6155));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6238), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6277));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6194), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6165), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6451));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6205), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6442), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6410), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6372));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6388), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6173), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6318));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6330), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6469), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6395));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6253), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6446), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6178));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I735 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6303), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6292));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20]));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5440));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[47]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6236));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6202));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6360));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6397));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6154), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6408));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I750 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6460), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I751 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6286), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I752 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6316), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6329), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6244));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6426), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6357));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6210), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6263), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6466));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6402), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6251));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6023));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5547));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I758 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[48]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[23]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I761 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I762 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6347));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6172));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6215));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6298), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6308), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6227));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I768 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6274), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6429), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I770 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6456), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6471), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6384));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I771 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6242), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6168));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6354), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6335), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6280));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I773 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6288), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6391));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I774 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[49]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5360), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5407));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[49]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6192));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6161));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I779 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6317));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I780 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6359));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I782 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6441), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6450), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6371));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I783 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6416), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6272), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6245), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6200));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6270), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6284), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6199));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6382), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6314));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6166), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6403), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6423));
XNOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6207));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I789 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10745));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6305));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6457));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6170));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6340));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I794 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I795 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6258), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6266), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6182));
OAI2BB2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I796 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6376), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6233), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6159), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6386));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I797 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6413), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6428), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6344));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I798 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6197), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6454));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6311), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6248), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6239));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6352));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25]));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I804 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6156), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6229));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I805 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6162), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6415), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6418));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6208));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I807 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6348), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6346), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6275));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I808 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6342), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6411));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I809 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6464), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6449));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I810 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I811 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6443), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6185));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I812 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6448), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6220), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6377));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I813 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6440), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6351));
OA21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I814 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6307), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6160), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6234));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I815 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I816 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6302), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6373));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I817 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6278), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6414), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6226));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I818 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I819 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I820 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6362), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6430));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I821 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6204));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I822 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6369), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6461), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6296));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I823 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6478), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6232), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6404));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I824 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6315), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6188));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I825 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I826 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17752));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I827 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6225), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6320), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6480));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I828 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17776));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I829 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6218), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6287));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I830 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17767), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17754), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17746));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I831 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I832 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6401), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6473));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6406), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6174), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6338));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6214), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6447));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6264), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6363), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6191));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6261), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6331));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6421), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6187), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6328));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I840 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779));
NOR2BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663));
NAND2BX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6763), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6839), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6779), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6764));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I848 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[3]));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I851 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I852 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7345));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I853 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7199));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6810));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I856 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6838), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I857 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I858 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6773), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6811), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6831));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I859 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6782), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6851));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I860 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620));
CLKINVX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I861 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I862 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I863 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I864 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I865 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7216));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I866 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I867 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7236));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I868 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I869 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I870 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I871 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I872 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6807), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6826));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6836), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6856));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6829), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6848), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6783));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6768), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6785), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6772));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6769), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6790));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6798), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6819));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6762), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6812), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6840));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I885 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6827), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6849));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I889 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6760));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[25]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10869));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6793), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6775), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6804));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I892 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6815), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6855));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I893 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6801), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6843));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I894 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[0]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I895 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I896 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I897 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7273));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I898 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I899 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I900 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I901 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I902 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17644));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I905 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7331));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I906 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7319), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I907 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I908 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6774), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6794));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6802), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6821));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6832), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6852));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I911 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6787));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6765), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6777), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6797));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6795), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6816));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I914 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6845));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I915 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6823), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6806), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6825));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I916 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6830), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6818), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6847));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6834), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6800));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I918 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1]));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I920 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I921 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7276), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7312), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[7]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I923 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I924 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I925 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7238), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I927 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I928 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I929 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I930 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7359), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10735), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I933 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7265), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I935 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7310), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I936 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7333), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7200), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I937 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7346), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I938 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I939 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I942 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7287), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7297), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I945 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7274), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I948 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7214), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7261), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7237), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I951 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I954 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7235), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10733));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I957 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I958 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I959 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7308), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I960 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I961 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7330), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I962 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7354), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7224), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I963 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7198), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I964 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7781), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7735), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I967 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I968 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7357), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7323), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7225), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7263), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7360), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7298), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I974 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7197));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I976 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I977 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10721), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10715));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I978 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7252), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I979 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7246), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I980 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I981 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10736), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[5]));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I982 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17664), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17618), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I983 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17637));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I984 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17974));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I985 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17642), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I986 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I987 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I988 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17660), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I989 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17628), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17638), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17663));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I990 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17653));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I991 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17626));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I992 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17620), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17632), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17649));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I993 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17631), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17648));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I994 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I995 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I996 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7253), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7290), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I997 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7348), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7218), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I998 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I999 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1000 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7289), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7215), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1001 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7324), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7251), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1002 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1003 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7705), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1004 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1005 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7335), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7229), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1006 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7202), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1007 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7326), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1008 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7361), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1009 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1010 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7242), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7267), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1011 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10737));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1012 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7284), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17655), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1013 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7219), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7240), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1014 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7363), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1015 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7230), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1016 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1017 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1018 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7316), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7304), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1019 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7255), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7277), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1020 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7232), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1021 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7266), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1022 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[23]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1023 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7221), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7340), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1024 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7292), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7313), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1025 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7269), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1026 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7209), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7303), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1027 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7798), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7688), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1028 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742), .AN(N7024), .B(N7088), .C(N7104));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1029 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7211));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1030 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7329), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1031 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7317), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1032 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7295), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1033 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7257), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1034 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7282), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1035 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7258), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1036 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1037 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7351));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1038 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7207), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1039 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7222), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1040 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7279));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1041 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7301), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1042 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7352), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1043 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4]));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5047 (.Y(N7928), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I5048 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800), .A(N7928));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1045 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7204));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1046 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7228), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1047 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7315), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1048 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558), .A(rm[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1049 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581), .A(rm[0]));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1050 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1051 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582), .A(rm[2]));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1052 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5), .A(rm[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1053 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1054 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48), .A(a_sign), .B(b_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4309));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1055 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1056 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6), .A(rm[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1057 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1058 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1059 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7322));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1060 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7280), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1061 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1062 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5955));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1063 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[24]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1064 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1065 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N626));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1066 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7524), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N627));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1067 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5967), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7503), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7530), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1068 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1069 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7336), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7603));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1070 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7606), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N1693), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1]));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1071 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4581), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7558));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1072 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1073 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7244));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1074 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__43), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[1]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1075 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7640), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7625), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__53));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1076 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N634), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__54));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1077 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7647), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N639));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1078 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7661));
CLKAND2X3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1079 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1080 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[2]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1081 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10790));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1082 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1083 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7761), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7751));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1084 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7742), .B(N7567));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1085 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[24]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10738));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1086 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7294), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7208), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1087 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7327), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7349), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7286));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1088 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7305), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7342), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1089 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7247), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7341), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7260));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1090 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7670), .B(N6842));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1091 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317), .A(rm[0]), .B(rm[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4582));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7567), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48));
AOI211XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1093 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8339), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8317), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N652), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1094 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961), .A(a_exp[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1095 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N573));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1096 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10851));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1097 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1098 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7961), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N560), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1099 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950), .A(a_exp[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7950), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N559), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4643), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N556), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980), .A(a_exp[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7980), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N562), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945), .A(a_exp[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7945), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N563), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970), .A(a_exp[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N561), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8025));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8024));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976), .A(a_exp[1]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7976), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N557), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941), .A(a_exp[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7941), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7972), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N558), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7946));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8015), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8021), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[13]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[16]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[9]));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[11]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7792));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[20]));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[17]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7769), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[23]));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[22]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7754), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7737));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7721), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7759));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7797), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7768));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[6]));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[7]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[3]));
CLKAND2X3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7667), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525), .A(N7646), .B(N6918));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17979));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23]), .A1(N7236), .B0(N7232));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62), .A(N7209), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N642));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .A(N6973), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317), .A(a_exp[0]), .B(a_exp[1]), .C(a_exp[7]), .D(a_exp[6]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4317), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4321));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354), .A(a_man[8]), .B(a_man[7]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352), .A(a_man[6]), .B(a_man[4]), .C(a_man[5]), .D(a_man[3]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4354), .B(a_man[10]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4352), .D(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377), .A(a_man[22]), .B(a_man[21]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4369), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4379));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340), .A(a_man[20]), .B(a_man[19]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1156 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4377), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4373), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4340));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1157 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338), .B(a_man[0]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10761), .D(a_man[1]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1158 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4357), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4346));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1159 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1160 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412), .A(b_exp[0]), .B(b_exp[1]), .C(b_exp[7]), .D(b_exp[6]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1161 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1162 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4412), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4416));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1163 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447), .A(b_man[6]), .B(b_man[4]), .C(b_man[5]), .D(b_man[3]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437), .A(b_man[10]), .B(b_man[8]), .C(b_man[9]), .D(b_man[7]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1166 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462), .A(b_man[0]), .B(b_man[1]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1167 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1168 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4464), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4474));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4433), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4462), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4468));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4447), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4437), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4454), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10769));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1172 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__15));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__10));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13));
AOI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1176 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[25]), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10775));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4525));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N7927));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1179 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8075), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7206), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[0]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1180 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[23]), .B(N7152));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1181 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513), .A(N7152), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17525));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17933), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17922));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8086), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8115), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8049));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513), .B(N7146));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[5]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8107));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8112), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8070));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8094), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8056));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1199 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7234), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1201 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10734), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[3]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1204 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7272), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__29[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7243));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8038), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8099));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087), .A0(N7251), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17513), .B0(N7249));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17529));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17517), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17541));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8071), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8088));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8045), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8109));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8106), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8083), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8078), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8066));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048), .A0(N7219), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076), .B0(N7217));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480), .A(N7138), .B(N7136), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17480), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8059), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2]), .A(N7184), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8090), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8110));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8067), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8084), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8055), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068), .A0(N7227), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8087), .B0(N7225));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5]), .A(N7178), .B(N7180), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8104), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8034));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8100), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8064));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8118), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8116), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8081));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3]), .A(N7192), .B(N7194), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8076));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8079), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8101));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8057), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8037), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8080), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7]), .A(N7170), .B(N7172), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8111), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8044), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8062));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6]), .A(N7162), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8082), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8053), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8072));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8068), .B(N7158));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4]));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17458), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17466), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17475));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6808), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6778));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17483), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17493), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8058), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8042), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8074));
OAI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489), .A0(N7203), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8048), .B0(N7199), .B1(N7201));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17489));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463), .A(N7051), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17456));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17485), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17470), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17463));
INVX6 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1255 (.Y(x[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8363), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7775), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7801), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7788));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7682), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7702));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7718), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7741));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7717), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7808), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704));
NAND4BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672), .AN(N7000), .B(N7070), .C(N7072), .D(N7074));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7757), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7772));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7732));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7804), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7748));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722), .A(N7575));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[21]), .A(N6835), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10843));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__13));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__18));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7025), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4931), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6802), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1273 (.Y(x[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8461), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7710), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7728), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7747));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7763), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7782));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7796), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7671));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7795), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7753), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786));
NAND4BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758), .AN(N7063), .B(N7079), .C(N7029), .D(N7083));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7693), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7708));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N2855));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7713), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689), .A(N7031));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7758), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[20]), .A(N6845), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10836));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4864), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6795), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1288 (.Y(x[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8435), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7686), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7724));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694), .AN(N7099), .B(N7095), .C(N7097));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7699));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7694), .B(N6933));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[19]), .A(N6855), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7679));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4796), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6722), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1297 (.Y(x[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8407), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7668), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7766), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7800));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773), .AN(N7039), .B(N7088), .C(N7090));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696), .A(N7642));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7773), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[18]), .A(N6850), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7731));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6984), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4884), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6715), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1306 (.Y(x[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8379), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7755), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7704), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7746));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803), .A(N7652));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829), .AN(N7006), .B(N7000), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676), .D(N7004));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[17]), .A(N6860), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10829));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7060), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4817), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6788), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1315 (.Y(x[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8353), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7691), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7786), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7678));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791), .AN(N7034), .B(N7063), .C(N7065));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7712));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7791), .B(N6997));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[16]), .A(N6819), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7684));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7000), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4901), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6708), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1324 (.Y(x[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8451), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7806), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7701), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7706));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[15]), .A(N6908), .B(N6910));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7076), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4839), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6701), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1330 (.Y(x[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8424), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716), .A(N7024), .B(N7567));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[14]), .A(N6868), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7716));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7016), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4922), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6694), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1336 (.Y(x[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8394), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822), .A(N7072), .B(N7575));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[13]), .A(N6913), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10822));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7092), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4854), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6781), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1342 (.Y(x[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8368), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815), .A(N7029), .B(N7031));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[12]), .A(N6888), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10815));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7035), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4791), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6774), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1348 (.Y(x[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8466), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10808), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7739), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7729));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[11]), .A(N6923), .B(N6925));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4875), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6767), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1354 (.Y(x[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8440), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801), .A(N7039), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[10]), .A(N6903), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10801));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7054), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4807), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6760), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1360 (.Y(x[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8412), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675), .A(N7006), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7803));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[9]), .A(N6878), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7675));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6995), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4893), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6687), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1366 (.Y(x[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8384), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794), .A(N7034), .B(N6997));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[8]), .A(N6893), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10794));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7071), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4829), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6753), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1372 (.Y(x[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8358), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[7]), .A(N6918), .B(N6920));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7011), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4912), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6680), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1377 (.Y(x[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8456), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[6]), .A(N7567), .B(N6900));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7086), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4847), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6746), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1382 (.Y(x[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8429), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7722), .B(N6885));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7028), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4934), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6673), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1387 (.Y(x[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8400), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[4]), .A(N6873), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7689));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6969), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4866), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6666), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1392 (.Y(x[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8373), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[3]), .A(N6933), .B(N6935));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7045), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4801), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6739), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1397 (.Y(x[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8346), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7696), .B(N6930));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6987), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4338), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6732), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1402 (.Y(x[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8445), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[1]), .A(N6938), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7676));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7064), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N4820), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6659), .S0(N7925));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1407 (.Y(x[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8417), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__55), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7776));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004), .A(b_man[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7004), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N5224), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__70), .B(N6725), .S0(N7927));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1412 (.Y(x[0]), .A(N6566), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8388), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8426));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8253), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__17), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .A(N6814), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__71));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1416 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1417 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1418 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1419 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1420 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1421 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[1]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1423 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8276), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8296), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
OR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N8243), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__8), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__4), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N635));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651), .A0(N6978), .A1(N6980), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__62));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[0]), .A(N6814), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1427 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N10742));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966), .A(a_sign), .B(b_sign));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N17966), .B0(a_sign), .B1(b_sign));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__16));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N645), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N6958));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7034), .B(b_sign));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017), .A(a_sign));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7050), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7096), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7017), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7090));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__6), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N706));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_1_I1438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[31]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7182), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7185), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_N7191));
EDFFHQX1 x_reg_31__I1470 (.Q(x[31]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[31]), .E(bdw_enable), .CK(aclk));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[0] = x[0];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[1] = x[1];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[2] = x[2];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[3] = x[3];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[4] = x[4];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[5] = x[5];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[6] = x[6];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[7] = x[7];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[8] = x[8];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[9] = x[9];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[10] = x[10];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[11] = x[11];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[12] = x[12];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[13] = x[13];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[14] = x[14];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[15] = x[15];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[16] = x[16];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[17] = x[17];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[18] = x[18];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[19] = x[19];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[20] = x[20];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[21] = x[21];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[22] = x[22];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[23] = x[23];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[24] = x[24];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[25] = x[25];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[26] = x[26];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[27] = x[27];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[28] = x[28];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[29] = x[29];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_x[30] = x[30];
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__27[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[30] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__35[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[34] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[35] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[38] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[39] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[40] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[43] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[44] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__50[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_0_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  vrPwTg/frhw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



