/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:24 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_4 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456;
wire N8516,N8554,N8561,N8568,N8574,N8577,N8586 
	,N8595,N8604,N8613,N8622,N8631,N8640,N8649,N8658 
	,N8667,N8676,N8685,N8694,N8703,N8712,N8721,N8730 
	,N8739,N8748,N8757,N8768,N8773,N8778,N8783,N8788 
	,N8793,N8798,N8803,N8808,N8813,N8818,N8823,N8828 
	,N8833,N8838,N8843,N8848,N8853,N8858,N8863,N8868 
	,N8873,N9105,N9131,N9157,N9493,N9495,N9532,N9534 
	,N9540,N9542,N9554,N9556,N9563,N9565,N9572,N9574 
	,N9581,N9583,N9600,N9602,N9609,N9611,N9618,N9620 
	,N9627,N9629,N9641,N9663,N9665,N9667,N9688,N9690 
	,N9695,N9711,N9713,N9715,N9836,N9838,N9846,N9848 
	,N9856,N9858,N9866,N9868,N9876,N9878,N9886,N9888 
	,N9942,N10007,N10009,N10017,N10019,N10064,N10066,N10076 
	,N10084,N10086,N10127,N10129,N10134,N10136,N10141,N10143 
	,N10148,N10155,N10157,N10164,N10171,N10176,N10178,N10183 
	,N10197,N10199,N10220,N10227,N10229,N10234,N10253,N10255 
	,N10931,N10932;
reg x_reg_21__retimed_I5715_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5715_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18];
	end
assign N10255 = x_reg_21__retimed_I5715_QOUT;
reg x_reg_21__retimed_I5714_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5714_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17];
	end
assign N10253 = x_reg_21__retimed_I5714_QOUT;
reg x_reg_21__retimed_I5706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5706_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19];
	end
assign N10234 = x_reg_21__retimed_I5706_QOUT;
reg x_reg_21__retimed_I5704_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5704_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21];
	end
assign N10229 = x_reg_21__retimed_I5704_QOUT;
reg x_reg_21__retimed_I5703_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5703_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20];
	end
assign N10227 = x_reg_21__retimed_I5703_QOUT;
reg x_reg_21__retimed_I5700_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5700_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0];
	end
assign N10220 = x_reg_21__retimed_I5700_QOUT;
reg x_reg_21__retimed_I5691_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5691_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16];
	end
assign N10199 = x_reg_21__retimed_I5691_QOUT;
reg x_reg_21__retimed_I5690_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5690_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15];
	end
assign N10197 = x_reg_21__retimed_I5690_QOUT;
reg x_reg_21__retimed_I5684_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5684_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3];
	end
assign N10183 = x_reg_21__retimed_I5684_QOUT;
reg x_reg_21__retimed_I5682_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5682_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12];
	end
assign N10178 = x_reg_21__retimed_I5682_QOUT;
reg x_reg_21__retimed_I5681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5681_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11];
	end
assign N10176 = x_reg_21__retimed_I5681_QOUT;
reg x_reg_21__retimed_I5679_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5679_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7];
	end
assign N10171 = x_reg_21__retimed_I5679_QOUT;
reg x_reg_21__retimed_I5676_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5676_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6];
	end
assign N10164 = x_reg_21__retimed_I5676_QOUT;
reg x_reg_21__retimed_I5673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5673_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14];
	end
assign N10157 = x_reg_21__retimed_I5673_QOUT;
reg x_reg_21__retimed_I5672_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5672_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13];
	end
assign N10155 = x_reg_21__retimed_I5672_QOUT;
reg x_reg_21__retimed_I5669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5669_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8];
	end
assign N10148 = x_reg_21__retimed_I5669_QOUT;
reg x_reg_21__retimed_I5667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5667_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2];
	end
assign N10143 = x_reg_21__retimed_I5667_QOUT;
reg x_reg_21__retimed_I5666_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5666_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1];
	end
assign N10141 = x_reg_21__retimed_I5666_QOUT;
reg x_reg_21__retimed_I5664_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5664_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10];
	end
assign N10136 = x_reg_21__retimed_I5664_QOUT;
reg x_reg_21__retimed_I5663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5663_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9];
	end
assign N10134 = x_reg_21__retimed_I5663_QOUT;
reg x_reg_21__retimed_I5661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5661_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5];
	end
assign N10129 = x_reg_21__retimed_I5661_QOUT;
reg x_reg_21__retimed_I5660_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5660_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4];
	end
assign N10127 = x_reg_21__retimed_I5660_QOUT;
reg x_reg_21__retimed_I5646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5646_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33];
	end
assign N10086 = x_reg_21__retimed_I5646_QOUT;
reg x_reg_21__retimed_I5645_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5645_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32];
	end
assign N10084 = x_reg_21__retimed_I5645_QOUT;
reg x_reg_21__retimed_I5643_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5643_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31];
	end
assign N10076 = x_reg_21__retimed_I5643_QOUT;
reg x_reg_21__retimed_I5640_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5640_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25];
	end
assign N10066 = x_reg_21__retimed_I5640_QOUT;
reg x_reg_21__retimed_I5639_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5639_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24];
	end
assign N10064 = x_reg_21__retimed_I5639_QOUT;
reg x_reg_21__retimed_I5623_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5623_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35];
	end
assign N10019 = x_reg_21__retimed_I5623_QOUT;
reg x_reg_21__retimed_I5622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5622_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34];
	end
assign N10017 = x_reg_21__retimed_I5622_QOUT;
reg x_reg_21__retimed_I5620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5620_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27];
	end
assign N10009 = x_reg_21__retimed_I5620_QOUT;
reg x_reg_21__retimed_I5619_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5619_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26];
	end
assign N10007 = x_reg_21__retimed_I5619_QOUT;
reg x_reg_21__retimed_I5595_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5595_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30];
	end
assign N9942 = x_reg_21__retimed_I5595_QOUT;
reg x_reg_21__retimed_I5577_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5577_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41];
	end
assign N9888 = x_reg_21__retimed_I5577_QOUT;
reg x_reg_21__retimed_I5576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5576_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40];
	end
assign N9886 = x_reg_21__retimed_I5576_QOUT;
reg x_reg_21__retimed_I5574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5574_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29];
	end
assign N9878 = x_reg_21__retimed_I5574_QOUT;
reg x_reg_21__retimed_I5573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5573_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28];
	end
assign N9876 = x_reg_21__retimed_I5573_QOUT;
reg x_reg_21__retimed_I5571_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5571_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45];
	end
assign N9868 = x_reg_21__retimed_I5571_QOUT;
reg x_reg_21__retimed_I5570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5570_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44];
	end
assign N9866 = x_reg_21__retimed_I5570_QOUT;
reg x_reg_21__retimed_I5568_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5568_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37];
	end
assign N9858 = x_reg_21__retimed_I5568_QOUT;
reg x_reg_21__retimed_I5567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5567_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36];
	end
assign N9856 = x_reg_21__retimed_I5567_QOUT;
reg x_reg_21__retimed_I5565_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5565_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39];
	end
assign N9848 = x_reg_21__retimed_I5565_QOUT;
reg x_reg_21__retimed_I5564_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5564_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38];
	end
assign N9846 = x_reg_21__retimed_I5564_QOUT;
reg x_reg_21__retimed_I5562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5562_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43];
	end
assign N9838 = x_reg_21__retimed_I5562_QOUT;
reg x_reg_21__retimed_I5561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5561_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42];
	end
assign N9836 = x_reg_21__retimed_I5561_QOUT;
reg x_reg_21__retimed_I5524_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5524_QOUT <= rm[2];
	end
assign N9715 = x_reg_21__retimed_I5524_QOUT;
reg x_reg_21__retimed_I5523_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5523_QOUT <= rm[0];
	end
assign N9713 = x_reg_21__retimed_I5523_QOUT;
reg x_reg_21__retimed_I5522_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5522_QOUT <= rm[1];
	end
assign N9711 = x_reg_21__retimed_I5522_QOUT;
reg x_reg_21__retimed_I5519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5519_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46];
	end
assign N9695 = x_reg_21__retimed_I5519_QOUT;
reg x_reg_21__retimed_I5517_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5517_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23];
	end
assign N9690 = x_reg_21__retimed_I5517_QOUT;
reg x_reg_21__retimed_I5516_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5516_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22];
	end
assign N9688 = x_reg_21__retimed_I5516_QOUT;
reg x_reg_21__retimed_I5507_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5507_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446;
	end
assign N9667 = x_reg_21__retimed_I5507_QOUT;
reg x_reg_21__retimed_I5506_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5506_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445;
	end
assign N9665 = x_reg_21__retimed_I5506_QOUT;
reg x_reg_21__retimed_I5505_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5505_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N9663 = x_reg_21__retimed_I5505_QOUT;
reg x_reg_21__retimed_I5497_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5497_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47];
	end
assign N9641 = x_reg_21__retimed_I5497_QOUT;
reg x_reg_21__retimed_I5496_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5496_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3];
	end
assign N9629 = x_reg_21__retimed_I5496_QOUT;
reg x_reg_21__retimed_I5495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5495_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3];
	end
assign N9627 = x_reg_21__retimed_I5495_QOUT;
reg x_reg_21__retimed_I5493_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5493_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
	end
assign N9620 = x_reg_21__retimed_I5493_QOUT;
reg x_reg_21__retimed_I5492_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5492_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7];
	end
assign N9618 = x_reg_21__retimed_I5492_QOUT;
reg x_reg_21__retimed_I5490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5490_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4];
	end
assign N9611 = x_reg_21__retimed_I5490_QOUT;
reg x_reg_21__retimed_I5489_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5489_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4];
	end
assign N9609 = x_reg_21__retimed_I5489_QOUT;
reg x_reg_21__retimed_I5487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5487_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2];
	end
assign N9602 = x_reg_21__retimed_I5487_QOUT;
reg x_reg_21__retimed_I5486_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5486_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2];
	end
assign N9600 = x_reg_21__retimed_I5486_QOUT;
reg x_reg_21__retimed_I5480_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5480_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1];
	end
assign N9583 = x_reg_21__retimed_I5480_QOUT;
reg x_reg_21__retimed_I5479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5479_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1];
	end
assign N9581 = x_reg_21__retimed_I5479_QOUT;
reg x_reg_21__retimed_I5477_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5477_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6];
	end
assign N9574 = x_reg_21__retimed_I5477_QOUT;
reg x_reg_21__retimed_I5476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5476_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6];
	end
assign N9572 = x_reg_21__retimed_I5476_QOUT;
reg x_reg_21__retimed_I5474_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5474_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5];
	end
assign N9565 = x_reg_21__retimed_I5474_QOUT;
reg x_reg_21__retimed_I5473_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5473_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5];
	end
assign N9563 = x_reg_21__retimed_I5473_QOUT;
reg x_reg_21__retimed_I5471_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5471_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0];
	end
assign N9556 = x_reg_21__retimed_I5471_QOUT;
reg x_reg_21__retimed_I5470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5470_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0];
	end
assign N9554 = x_reg_21__retimed_I5470_QOUT;
reg x_reg_21__retimed_I5466_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5466_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8];
	end
assign N9542 = x_reg_21__retimed_I5466_QOUT;
reg x_reg_21__retimed_I5465_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5465_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8];
	end
assign N9540 = x_reg_21__retimed_I5465_QOUT;
reg x_reg_21__retimed_I5463_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5463_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9];
	end
assign N9534 = x_reg_21__retimed_I5463_QOUT;
reg x_reg_21__retimed_I5462_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5462_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9];
	end
assign N9532 = x_reg_21__retimed_I5462_QOUT;
reg x_reg_21__retimed_I5447_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5447_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27;
	end
assign N9495 = x_reg_21__retimed_I5447_QOUT;
reg x_reg_21__retimed_I5446_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5446_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
	end
assign N9493 = x_reg_21__retimed_I5446_QOUT;
reg x_reg_21__retimed_I5331_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5331_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26;
	end
assign N9157 = x_reg_21__retimed_I5331_QOUT;
reg x_reg_21__retimed_I5329_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5329_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144;
	end
assign N9131 = x_reg_21__retimed_I5329_QOUT;
reg x_reg_21__retimed_I5327_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5327_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225;
	end
assign N9105 = x_reg_21__retimed_I5327_QOUT;
reg x_reg_21__retimed_I5234_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5234_QOUT <= a_man[21];
	end
assign N8873 = x_reg_21__retimed_I5234_QOUT;
reg x_reg_20__retimed_I5232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I5232_QOUT <= a_man[20];
	end
assign N8868 = x_reg_20__retimed_I5232_QOUT;
reg x_reg_19__retimed_I5230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I5230_QOUT <= a_man[19];
	end
assign N8863 = x_reg_19__retimed_I5230_QOUT;
reg x_reg_18__retimed_I5228_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I5228_QOUT <= a_man[18];
	end
assign N8858 = x_reg_18__retimed_I5228_QOUT;
reg x_reg_17__retimed_I5226_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I5226_QOUT <= a_man[17];
	end
assign N8853 = x_reg_17__retimed_I5226_QOUT;
reg x_reg_16__retimed_I5224_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I5224_QOUT <= a_man[16];
	end
assign N8848 = x_reg_16__retimed_I5224_QOUT;
reg x_reg_15__retimed_I5222_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I5222_QOUT <= a_man[15];
	end
assign N8843 = x_reg_15__retimed_I5222_QOUT;
reg x_reg_14__retimed_I5220_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I5220_QOUT <= a_man[14];
	end
assign N8838 = x_reg_14__retimed_I5220_QOUT;
reg x_reg_13__retimed_I5218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I5218_QOUT <= a_man[13];
	end
assign N8833 = x_reg_13__retimed_I5218_QOUT;
reg x_reg_12__retimed_I5216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I5216_QOUT <= a_man[12];
	end
assign N8828 = x_reg_12__retimed_I5216_QOUT;
reg x_reg_11__retimed_I5214_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I5214_QOUT <= a_man[11];
	end
assign N8823 = x_reg_11__retimed_I5214_QOUT;
reg x_reg_10__retimed_I5212_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I5212_QOUT <= a_man[10];
	end
assign N8818 = x_reg_10__retimed_I5212_QOUT;
reg x_reg_9__retimed_I5210_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I5210_QOUT <= a_man[9];
	end
assign N8813 = x_reg_9__retimed_I5210_QOUT;
reg x_reg_8__retimed_I5208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I5208_QOUT <= a_man[8];
	end
assign N8808 = x_reg_8__retimed_I5208_QOUT;
reg x_reg_7__retimed_I5206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I5206_QOUT <= a_man[7];
	end
assign N8803 = x_reg_7__retimed_I5206_QOUT;
reg x_reg_6__retimed_I5204_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I5204_QOUT <= a_man[6];
	end
assign N8798 = x_reg_6__retimed_I5204_QOUT;
reg x_reg_5__retimed_I5202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I5202_QOUT <= a_man[5];
	end
assign N8793 = x_reg_5__retimed_I5202_QOUT;
reg x_reg_4__retimed_I5200_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I5200_QOUT <= a_man[4];
	end
assign N8788 = x_reg_4__retimed_I5200_QOUT;
reg x_reg_3__retimed_I5198_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I5198_QOUT <= a_man[3];
	end
assign N8783 = x_reg_3__retimed_I5198_QOUT;
reg x_reg_2__retimed_I5196_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I5196_QOUT <= a_man[2];
	end
assign N8778 = x_reg_2__retimed_I5196_QOUT;
reg x_reg_1__retimed_I5194_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I5194_QOUT <= a_man[1];
	end
assign N8773 = x_reg_1__retimed_I5194_QOUT;
reg x_reg_0__retimed_I5192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I5192_QOUT <= a_man[0];
	end
assign N8768 = x_reg_0__retimed_I5192_QOUT;
reg x_reg_21__retimed_I5187_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I5187_QOUT <= b_man[21];
	end
assign N8757 = x_reg_21__retimed_I5187_QOUT;
reg x_reg_20__retimed_I5183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I5183_QOUT <= b_man[20];
	end
assign N8748 = x_reg_20__retimed_I5183_QOUT;
reg x_reg_19__retimed_I5179_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I5179_QOUT <= b_man[19];
	end
assign N8739 = x_reg_19__retimed_I5179_QOUT;
reg x_reg_18__retimed_I5175_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I5175_QOUT <= b_man[18];
	end
assign N8730 = x_reg_18__retimed_I5175_QOUT;
reg x_reg_17__retimed_I5171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I5171_QOUT <= b_man[17];
	end
assign N8721 = x_reg_17__retimed_I5171_QOUT;
reg x_reg_16__retimed_I5167_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I5167_QOUT <= b_man[16];
	end
assign N8712 = x_reg_16__retimed_I5167_QOUT;
reg x_reg_15__retimed_I5163_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I5163_QOUT <= b_man[15];
	end
assign N8703 = x_reg_15__retimed_I5163_QOUT;
reg x_reg_14__retimed_I5159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I5159_QOUT <= b_man[14];
	end
assign N8694 = x_reg_14__retimed_I5159_QOUT;
reg x_reg_13__retimed_I5155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I5155_QOUT <= b_man[13];
	end
assign N8685 = x_reg_13__retimed_I5155_QOUT;
reg x_reg_12__retimed_I5151_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I5151_QOUT <= b_man[12];
	end
assign N8676 = x_reg_12__retimed_I5151_QOUT;
reg x_reg_11__retimed_I5147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I5147_QOUT <= b_man[11];
	end
assign N8667 = x_reg_11__retimed_I5147_QOUT;
reg x_reg_10__retimed_I5143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I5143_QOUT <= b_man[10];
	end
assign N8658 = x_reg_10__retimed_I5143_QOUT;
reg x_reg_9__retimed_I5139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I5139_QOUT <= b_man[9];
	end
assign N8649 = x_reg_9__retimed_I5139_QOUT;
reg x_reg_8__retimed_I5135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I5135_QOUT <= b_man[8];
	end
assign N8640 = x_reg_8__retimed_I5135_QOUT;
reg x_reg_7__retimed_I5131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I5131_QOUT <= b_man[7];
	end
assign N8631 = x_reg_7__retimed_I5131_QOUT;
reg x_reg_6__retimed_I5127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I5127_QOUT <= b_man[6];
	end
assign N8622 = x_reg_6__retimed_I5127_QOUT;
reg x_reg_5__retimed_I5123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I5123_QOUT <= b_man[5];
	end
assign N8613 = x_reg_5__retimed_I5123_QOUT;
reg x_reg_4__retimed_I5119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I5119_QOUT <= b_man[4];
	end
assign N8604 = x_reg_4__retimed_I5119_QOUT;
reg x_reg_3__retimed_I5115_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I5115_QOUT <= b_man[3];
	end
assign N8595 = x_reg_3__retimed_I5115_QOUT;
reg x_reg_2__retimed_I5111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I5111_QOUT <= b_man[2];
	end
assign N8586 = x_reg_2__retimed_I5111_QOUT;
reg x_reg_1__retimed_I5107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I5107_QOUT <= b_man[1];
	end
assign N8577 = x_reg_1__retimed_I5107_QOUT;
reg x_reg_0__retimed_I5106_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I5106_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
	end
assign N8574 = x_reg_0__retimed_I5106_QOUT;
assign N10931 = !N8574;
assign N10932 = !N10931;
reg x_reg_0__retimed_I5103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I5103_QOUT <= b_man[0];
	end
assign N8568 = x_reg_0__retimed_I5103_QOUT;
reg x_reg_22__retimed_I5100_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I5100_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055;
	end
assign N8561 = x_reg_22__retimed_I5100_QOUT;
reg x_reg_23__retimed_I5097_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I5097_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025;
	end
assign N8554 = x_reg_23__retimed_I5097_QOUT;
reg x_reg_29__retimed_I5081_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_29__retimed_I5081_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008;
	end
assign N8516 = x_reg_29__retimed_I5081_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007 = !(a_exp[0] & a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434 = !((a_exp[7] & a_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896 = !(b_exp[0] & b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426 = !((b_exp[7] & b_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936 = !(((b_man[0] | b_man[1]) | b_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919 = !(b_man[10] | b_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938 = !(b_man[6] | b_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927 = !(b_man[8] | b_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947 = !(b_man[4] | b_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092 = !(b_exp[0] | b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099 = !(b_exp[5] | b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096 = !(b_exp[7] | b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087 = !(b_exp[3] | b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0] = (!b_exp[0]) ^ a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318 = (!b_man[22]) ^ b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217 = !a_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504 = !a_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862 = !a_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011 = b_man[22] | b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392 = (!b_man[20]) ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007 = b_man[21] ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552 = !b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415 = !a_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152 = !a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716 = !a_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076 = !a_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169 = b_man[19] ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463 = (!b_man[18]) ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407 = !b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529 = (!b_man[16]) ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973 = b_man[17] ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268 = !b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616 = !a_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352 = !a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924 = !a_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276 = !a_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212 = !a_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566 = !a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124 = !b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598 = (!b_man[14]) ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751 = b_man[15] ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664 = (!b_man[12]) ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942 = b_man[13] ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981 = !b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720 = b_man[11] ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737 = (!b_man[10]) ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827 = !b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131 = !a_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473 = !a_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417 = !a_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779 = !a_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805 = (!b_man[8]) ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911 = b_man[9] ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678 = !b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334 = !a_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675 = !a_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871 = (!b_man[6]) ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691 = b_man[7] ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531 = !b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881 = b_man[5] ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941 = (!b_man[4]) ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377 = !b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624 = !a_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988 = !a_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014 = (!b_man[2]) ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662 = b_man[3] ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237 = !b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268 = !a_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357 = !b_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361 = !b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529 = !a_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831 = !(b_man[21] & b_man[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543 = !(b_man[19] & b_man[20]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901 = b_man[21] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610 = !(b_man[17] & b_man[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971 = b_man[19] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676 = !(b_man[15] & b_man[16]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043 = b_man[17] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749 = !(b_man[13] & b_man[14]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105 = b_man[15] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817 = !(b_man[11] & b_man[12]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172 = b_man[13] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883 = !(b_man[9] & b_man[10]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236 = b_man[11] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952 = !(b_man[7] & b_man[8]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301 = b_man[9] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028 = !(b_man[5] & b_man[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369 = b_man[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090 = !(b_man[3] & b_man[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430 = b_man[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154 = !(b_man[1] & b_man[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495 = b_man[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364) & (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513) | (!(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 = N9641;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 | N9695);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9866) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9838);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9838) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9836);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9695) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9868);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9868) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9866);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9856) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10019);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10019) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10017);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9846) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9858);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10017) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10086);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10086) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10084);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10084) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10076);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10076) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9942);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9858) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9856);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9876) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10009);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10009) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10007);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9942) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9878);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10007) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10066);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10066) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10064);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10064) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9690);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9878) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9876);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9836) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9888);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9888) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9886);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9886) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9848);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9848) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9846);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9690) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N9688);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23 = a_sign ^ b_sign;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10143) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10141);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10164) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10129);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10127) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10183);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10148) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10171);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10136) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10134);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10157) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10155);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10178) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10176);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10199) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10129) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10127);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10134) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10148);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10171) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10164);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10176) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10136);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10183) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10143);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N9688) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10229);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10227) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10234);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10255) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10253);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0] = b_man[1] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10220;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10141) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10220);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10229) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10227);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10155) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10178);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10253) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10199);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10197) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10157);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360 & N10234) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360) & N10255);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443) | N9711) | N9713) | N9715);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447 = ((N9663 | N9665) | N9667) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450 = ((!N9667) & (!N9665)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24]) | N9641);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9556) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9554);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765 = b_exp[0] | a_exp[0];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]} = {1'B0, a_exp[1]} + {1'B0, b_exp[1]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2]} = {1'B0, a_exp[2]} + {1'B0, b_exp[2]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9602) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9600);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3]} = {1'B0, a_exp[3]} + {1'B0, b_exp[3]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]} = {1'B0, a_exp[4]} + {1'B0, b_exp[4]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9611) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9609);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]} = {1'B0, a_exp[5]} + {1'B0, b_exp[5]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9565) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9563);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]} = {1'B0, a_exp[6]} + {1'B0, b_exp[6]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761 = !a_exp[7];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]} = {1'B0, b_exp[7]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9620) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9618);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9629) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9627);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] = (!a_exp[7]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9542) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9540);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9574) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9572);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9583) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9581);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9] = !(a_exp[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38 & N9534) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38) & N9532);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964 = !(((N9493 | N9495) | N9157) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 = !(N9105 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8873);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 = !(N9131 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 = !(N9157 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986 = !(rm[0] & rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7 = !(rm[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8757) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[21] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8868);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8748) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[20] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8863);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8739) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[19] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8858);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8730) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[18] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8853);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8721) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[17] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8848);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8712) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[16] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8843);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8703) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[15] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8838);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8694) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[14] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8833);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8685) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[13] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8828);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8676) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[12] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8823);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8667) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[11] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8818);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8658) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[10] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8813);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8649) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[9] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8808);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8640) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[8] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8803);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8631) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8798);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8622) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8793);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8613) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[5] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8788);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27] & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8604) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8783);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8595) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[3] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8778);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8586) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[2] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8773);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8577) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[1] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082 & N8768);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192 & N8568) | (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106 & N10932));
assign x[0] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47);
assign x[22] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8561) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008 = float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470;
assign x[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7]);
assign x[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]);
assign x[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]);
assign x[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]);
assign x[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]);
assign x[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]);
assign x[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8516) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004 = !float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42) | float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470);
assign x[23] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49 & N8554) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22 & (!b_sign));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136 = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15 & a_sign) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26) & float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23);
reg x_reg_31__I1669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__I1669_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31];
	end
assign x[31] = x_reg_31__I1669_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vrn1SgnYoxo= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



