/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:28 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_5 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456;
wire N4120,N8900,N8938,N8945,N8952,N8958,N8961 
	,N8970,N8979,N8988,N8997,N9006,N9015,N9024,N9033 
	,N9042,N9051,N9060,N9069,N9078,N9087,N9096,N9105 
	,N9114,N9123,N9132,N9141,N9152,N9157,N9162,N9167 
	,N9172,N9177,N9182,N9187,N9192,N9197,N9202,N9207 
	,N9212,N9217,N9222,N9227,N9232,N9237,N9242,N9247 
	,N9252,N9257,N9624,N9631,N9633,N9638,N9645,N9652 
	,N9659,N9666,N9671,N9673,N9678,N9680,N9706,N9732 
	,N9758,N9925,N9931,N9934,N9943,N9952,N9961,N9970 
	,N9979,N9988,N9997,N10006,N10015,N10024,N10033,N10042 
	,N10051,N10060,N10069,N10078,N10087,N10096,N10105,N10114 
	,N10125,N10130,N10135,N10140,N10145,N10150,N10155,N10160 
	,N10165,N10170,N10175,N10180,N10185,N10190,N10195,N10200 
	,N10205,N10210,N10215,N10220,N10225,N10230,N10233,N10239 
	,N10242,N10248,N10251,N10257,N10260,N10266,N10269,N10275 
	,N10278,N10284,N10287,N10293,N10296,N10302,N10305,N10311 
	,N10314,N10320,N10323,N10329,N10332,N10338,N10341,N10347 
	,N10350,N10356,N10359,N10365,N10368,N10374,N10377,N10383 
	,N10386,N10392,N10395,N10401,N10404,N10410,N10413,N10419 
	,N10422,N10428,N10567,N10593,N10619,N10645,N10751,N10753 
	,N10790,N10792,N10798,N10800,N10812,N10814,N10821,N10823 
	,N10830,N10832,N10839,N10841,N10858,N10860,N10867,N10869 
	,N10876,N10878,N10885,N10887,N10921,N10923,N10925,N10969 
	,N10971,N10973,N11301,N11307,N11313,N11319,N11325,N11331 
	,N11337,N11343,N11349,N11355,N11361,N11451,N11453,N11458 
	,N11460,N11465,N11467,N11472,N11479,N11481,N11488,N11495 
	,N11500,N11502,N11507,N11521,N11523,N11536,N11539,N11549 
	,N11552,N11559,N11566,N11573,N11583,N11589,N11592,N11610 
	,N11624,N11643,N11645,N11658,N11662,N11664,N11672,N11678 
	,N11684,N11692,N11694,N11702,N11710,N11712,N11717,N11727 
	,N11733,N11739,N11742,N11752,N11756,N11758,N11791,N11793 
	,N11802,N11804,N11810,N11812,N11821,N11823,N11829,N11831 
	,N11835,N11837,N11840,N11904,N11906,N11930,N11941,N11949 
	,N11951,N11960,N11962,N11971,N11973,N11981,N11983,N12644 
	,N12649,N12652,N12655,N12658,N12662,N13247,N13248,N13249 
	,N13250,N13251,N13252,N13253,N13254,N13255,N13256,N13257 
	,N13258,N13259,N13260,N13261,N13262,N13263,N13264,N13265 
	,N13266,N13267,N13268,N13270,N13271,N13273,N13280,N13287 
	,N13294,N13303,N13309,N13311,N13319;
reg x_reg_L1_21__retimed_I6582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6582_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49;
	end
assign N12662 = x_reg_L1_21__retimed_I6582_QOUT;
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6870 (.Y(N13247), .A(N12662));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6871 (.Y(N13248), .A(N13247));
reg x_reg_L0_21__retimed_I6580_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6580_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384;
	end
assign N12658 = x_reg_L0_21__retimed_I6580_QOUT;
reg x_reg_L0_21__retimed_I6579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6579_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751;
	end
assign N12655 = x_reg_L0_21__retimed_I6579_QOUT;
reg x_reg_L0_21__retimed_I6578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6578_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275;
	end
assign N12652 = x_reg_L0_21__retimed_I6578_QOUT;
reg x_reg_L0_21__retimed_I6577_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6577_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613;
	end
assign N12649 = x_reg_L0_21__retimed_I6577_QOUT;
reg x_reg_L0_21__retimed_I6575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6575_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20];
	end
assign N12644 = x_reg_L0_21__retimed_I6575_QOUT;
reg x_reg_L0_21__retimed_I6291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6291_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922;
	end
assign N11983 = x_reg_L0_21__retimed_I6291_QOUT;
reg x_reg_L0_21__retimed_I6290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6290_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563;
	end
assign N11981 = x_reg_L0_21__retimed_I6290_QOUT;
reg x_reg_L0_21__retimed_I6288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6288_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016;
	end
assign N11973 = x_reg_L0_21__retimed_I6288_QOUT;
reg x_reg_L0_21__retimed_I6287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6287_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651;
	end
assign N11971 = x_reg_L0_21__retimed_I6287_QOUT;
reg x_reg_L0_21__retimed_I6284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6284_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501;
	end
assign N11962 = x_reg_L0_21__retimed_I6284_QOUT;
reg x_reg_L0_21__retimed_I6283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6283_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099;
	end
assign N11960 = x_reg_L0_21__retimed_I6283_QOUT;
reg x_reg_L0_21__retimed_I6280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6280_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415;
	end
assign N11951 = x_reg_L0_21__retimed_I6280_QOUT;
reg x_reg_L0_21__retimed_I6279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6279_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342;
	end
assign N11949 = x_reg_L0_21__retimed_I6279_QOUT;
reg x_reg_L0_21__retimed_I6276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6276_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811;
	end
assign N11941 = x_reg_L0_21__retimed_I6276_QOUT;
reg x_reg_L0_21__retimed_I6272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6272_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244;
	end
assign N11930 = x_reg_L0_21__retimed_I6272_QOUT;
reg x_reg_L0_21__retimed_I6264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6264_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824;
	end
assign N11906 = x_reg_L0_21__retimed_I6264_QOUT;
reg x_reg_L0_21__retimed_I6263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6263_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185;
	end
assign N11904 = x_reg_L0_21__retimed_I6263_QOUT;
reg x_reg_L0_21__retimed_I6257_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6257_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656;
	end
assign N11840 = x_reg_L0_21__retimed_I6257_QOUT;
reg x_reg_L0_21__retimed_I6256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6256_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314;
	end
assign N11837 = x_reg_L0_21__retimed_I6256_QOUT;
reg x_reg_L0_21__retimed_I6255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6255_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495;
	end
assign N11835 = x_reg_L0_21__retimed_I6255_QOUT;
reg x_reg_L0_21__retimed_I6254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6254_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396;
	end
assign N11831 = x_reg_L0_21__retimed_I6254_QOUT;
reg x_reg_L0_21__retimed_I6253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6253_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471;
	end
assign N11829 = x_reg_L0_21__retimed_I6253_QOUT;
reg x_reg_L0_21__retimed_I6251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6251_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694;
	end
assign N11823 = x_reg_L0_21__retimed_I6251_QOUT;
reg x_reg_L0_21__retimed_I6250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6250_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435;
	end
assign N11821 = x_reg_L0_21__retimed_I6250_QOUT;
reg x_reg_L0_21__retimed_I6247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6247_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413;
	end
assign N11812 = x_reg_L0_21__retimed_I6247_QOUT;
reg x_reg_L0_21__retimed_I6246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6246_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073;
	end
assign N11810 = x_reg_L0_21__retimed_I6246_QOUT;
reg x_reg_L0_21__retimed_I6244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6244_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171;
	end
assign N11804 = x_reg_L0_21__retimed_I6244_QOUT;
reg x_reg_L0_21__retimed_I6243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6243_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524;
	end
assign N11802 = x_reg_L0_21__retimed_I6243_QOUT;
reg x_reg_L0_21__retimed_I6240_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6240_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669;
	end
assign N11793 = x_reg_L0_21__retimed_I6240_QOUT;
reg x_reg_L0_21__retimed_I6239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6239_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036;
	end
assign N11791 = x_reg_L0_21__retimed_I6239_QOUT;
reg x_reg_L0_21__retimed_I6225_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6225_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539;
	end
assign N11758 = x_reg_L0_21__retimed_I6225_QOUT;
reg x_reg_L0_21__retimed_I6224_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6224_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185;
	end
assign N11756 = x_reg_L0_21__retimed_I6224_QOUT;
reg x_reg_L0_21__retimed_I6223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6223_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112;
	end
assign N11752 = x_reg_L0_21__retimed_I6223_QOUT;
reg x_reg_L0_21__retimed_I6219_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6219_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256;
	end
assign N11742 = x_reg_L0_21__retimed_I6219_QOUT;
reg x_reg_L0_21__retimed_I6218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6218_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193;
	end
assign N11739 = x_reg_L0_21__retimed_I6218_QOUT;
reg x_reg_L0_21__retimed_I6216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6216_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904;
	end
assign N11733 = x_reg_L0_21__retimed_I6216_QOUT;
reg x_reg_L0_21__retimed_I6214_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6214_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596;
	end
assign N11727 = x_reg_L0_21__retimed_I6214_QOUT;
reg x_reg_L0_21__retimed_I6210_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6210_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423;
	end
assign N11717 = x_reg_L0_21__retimed_I6210_QOUT;
reg x_reg_L0_21__retimed_I6208_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6208_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733;
	end
assign N11712 = x_reg_L0_21__retimed_I6208_QOUT;
reg x_reg_L0_21__retimed_I6207_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6207_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389;
	end
assign N11710 = x_reg_L0_21__retimed_I6207_QOUT;
reg x_reg_L0_21__retimed_I6205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6205_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197;
	end
assign N11702 = x_reg_L0_21__retimed_I6205_QOUT;
reg x_reg_L0_21__retimed_I6202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6202_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527;
	end
assign N11694 = x_reg_L0_21__retimed_I6202_QOUT;
reg x_reg_L0_21__retimed_I6201_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6201_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191;
	end
assign N11692 = x_reg_L0_21__retimed_I6201_QOUT;
reg x_reg_L0_21__retimed_I6199_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6199_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787;
	end
assign N11684 = x_reg_L0_21__retimed_I6199_QOUT;
reg x_reg_L0_21__retimed_I6197_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6197_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274;
	end
assign N11678 = x_reg_L0_21__retimed_I6197_QOUT;
reg x_reg_L0_21__retimed_I6195_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6195_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995;
	end
assign N11672 = x_reg_L0_21__retimed_I6195_QOUT;
reg x_reg_L0_21__retimed_I6192_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6192_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333;
	end
assign N11664 = x_reg_L0_21__retimed_I6192_QOUT;
reg x_reg_L0_21__retimed_I6191_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6191_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986;
	end
assign N11662 = x_reg_L0_21__retimed_I6191_QOUT;
reg x_reg_L0_21__retimed_I6190_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6190_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680;
	end
assign N11658 = x_reg_L0_21__retimed_I6190_QOUT;
reg x_reg_L0_21__retimed_I6185_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6185_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18];
	end
assign N11645 = x_reg_L0_21__retimed_I6185_QOUT;
reg x_reg_L0_21__retimed_I6184_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6184_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17];
	end
assign N11643 = x_reg_L0_21__retimed_I6184_QOUT;
reg x_reg_L0_21__retimed_I6176_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6176_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19];
	end
assign N11624 = x_reg_L0_21__retimed_I6176_QOUT;
reg x_reg_L0_21__retimed_I6170_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6170_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0];
	end
assign N11610 = x_reg_L0_21__retimed_I6170_QOUT;
reg x_reg_L0_21__retimed_I6162_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6162_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055;
	end
assign N11592 = x_reg_L0_21__retimed_I6162_QOUT;
reg x_reg_L0_21__retimed_I6161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6161_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395;
	end
assign N11589 = x_reg_L0_21__retimed_I6161_QOUT;
reg x_reg_L0_21__retimed_I6159_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6159_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692;
	end
assign N11583 = x_reg_L0_21__retimed_I6159_QOUT;
reg x_reg_L0_21__retimed_I6155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6155_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219;
	end
assign N11573 = x_reg_L0_21__retimed_I6155_QOUT;
reg x_reg_L0_21__retimed_I6152_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6152_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623;
	end
assign N11566 = x_reg_L0_21__retimed_I6152_QOUT;
reg x_reg_L0_21__retimed_I6149_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6149_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422;
	end
assign N11559 = x_reg_L0_21__retimed_I6149_QOUT;
reg x_reg_L0_21__retimed_I6146_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6146_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225;
	end
assign N11552 = x_reg_L0_21__retimed_I6146_QOUT;
reg x_reg_L0_21__retimed_I6145_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6145_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571;
	end
assign N11549 = x_reg_L0_21__retimed_I6145_QOUT;
reg x_reg_L0_21__retimed_I6141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6141_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025;
	end
assign N11539 = x_reg_L0_21__retimed_I6141_QOUT;
reg x_reg_L0_21__retimed_I6140_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6140_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480;
	end
assign N11536 = x_reg_L0_21__retimed_I6140_QOUT;
reg x_reg_L0_21__retimed_I6135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6135_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16];
	end
assign N11523 = x_reg_L0_21__retimed_I6135_QOUT;
reg x_reg_L0_21__retimed_I6134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6134_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15];
	end
assign N11521 = x_reg_L0_21__retimed_I6134_QOUT;
reg x_reg_L0_21__retimed_I6128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6128_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3];
	end
assign N11507 = x_reg_L0_21__retimed_I6128_QOUT;
reg x_reg_L0_21__retimed_I6126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6126_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12];
	end
assign N11502 = x_reg_L0_21__retimed_I6126_QOUT;
reg x_reg_L0_21__retimed_I6125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6125_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11];
	end
assign N11500 = x_reg_L0_21__retimed_I6125_QOUT;
reg x_reg_L0_21__retimed_I6123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6123_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7];
	end
assign N11495 = x_reg_L0_21__retimed_I6123_QOUT;
reg x_reg_L0_21__retimed_I6120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6120_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6];
	end
assign N11488 = x_reg_L0_21__retimed_I6120_QOUT;
reg x_reg_L0_21__retimed_I6117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6117_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14];
	end
assign N11481 = x_reg_L0_21__retimed_I6117_QOUT;
reg x_reg_L0_21__retimed_I6116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6116_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13];
	end
assign N11479 = x_reg_L0_21__retimed_I6116_QOUT;
reg x_reg_L0_21__retimed_I6113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6113_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8];
	end
assign N11472 = x_reg_L0_21__retimed_I6113_QOUT;
reg x_reg_L0_21__retimed_I6111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6111_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2];
	end
assign N11467 = x_reg_L0_21__retimed_I6111_QOUT;
reg x_reg_L0_21__retimed_I6110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6110_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1];
	end
assign N11465 = x_reg_L0_21__retimed_I6110_QOUT;
reg x_reg_L0_21__retimed_I6108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6108_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10];
	end
assign N11460 = x_reg_L0_21__retimed_I6108_QOUT;
reg x_reg_L0_21__retimed_I6107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6107_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9];
	end
assign N11458 = x_reg_L0_21__retimed_I6107_QOUT;
reg x_reg_L0_21__retimed_I6105_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6105_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5];
	end
assign N11453 = x_reg_L0_21__retimed_I6105_QOUT;
reg x_reg_L0_21__retimed_I6104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6104_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4];
	end
assign N11451 = x_reg_L0_21__retimed_I6104_QOUT;
reg x_reg_L0_21__retimed_I6073_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6073_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483;
	end
assign N11361 = x_reg_L0_21__retimed_I6073_QOUT;
reg x_reg_L0_21__retimed_I6071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6071_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360;
	end
assign N11355 = x_reg_L0_21__retimed_I6071_QOUT;
reg x_reg_L0_21__retimed_I6069_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6069_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161;
	end
assign N11349 = x_reg_L0_21__retimed_I6069_QOUT;
reg x_reg_L0_21__retimed_I6067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6067_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564;
	end
assign N11343 = x_reg_L0_21__retimed_I6067_QOUT;
reg x_reg_L0_21__retimed_I6065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6065_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284;
	end
assign N11337 = x_reg_L0_21__retimed_I6065_QOUT;
reg x_reg_L0_21__retimed_I6063_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6063_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082;
	end
assign N11331 = x_reg_L0_21__retimed_I6063_QOUT;
reg x_reg_L0_21__retimed_I6061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6061_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367;
	end
assign N11325 = x_reg_L0_21__retimed_I6061_QOUT;
reg x_reg_L0_21__retimed_I6059_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6059_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166;
	end
assign N11319 = x_reg_L0_21__retimed_I6059_QOUT;
reg x_reg_L0_21__retimed_I6057_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6057_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869;
	end
assign N11313 = x_reg_L0_21__retimed_I6057_QOUT;
reg x_reg_L0_21__retimed_I6055_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6055_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659;
	end
assign N11307 = x_reg_L0_21__retimed_I6055_QOUT;
reg x_reg_L0_21__retimed_I6053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6053_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449;
	end
assign N11301 = x_reg_L0_21__retimed_I6053_QOUT;
reg x_reg_L0_21__retimed_I5946_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5946_QOUT <= rm[2];
	end
assign N10973 = x_reg_L0_21__retimed_I5946_QOUT;
reg x_reg_L0_21__retimed_I5945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5945_QOUT <= rm[0];
	end
assign N10971 = x_reg_L0_21__retimed_I5945_QOUT;
reg x_reg_L0_21__retimed_I5944_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5944_QOUT <= rm[1];
	end
assign N10969 = x_reg_L0_21__retimed_I5944_QOUT;
reg x_reg_L0_21__retimed_I5929_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5929_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446;
	end
assign N10925 = x_reg_L0_21__retimed_I5929_QOUT;
reg x_reg_L0_21__retimed_I5928_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5928_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445;
	end
assign N10923 = x_reg_L0_21__retimed_I5928_QOUT;
reg x_reg_L0_21__retimed_I5927_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5927_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N10921 = x_reg_L0_21__retimed_I5927_QOUT;
reg x_reg_L0_21__retimed_I5918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5918_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3];
	end
assign N10887 = x_reg_L0_21__retimed_I5918_QOUT;
reg x_reg_L0_21__retimed_I5917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5917_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3];
	end
assign N10885 = x_reg_L0_21__retimed_I5917_QOUT;
reg x_reg_L0_21__retimed_I5915_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5915_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7];
	end
assign N10878 = x_reg_L0_21__retimed_I5915_QOUT;
reg x_reg_L0_21__retimed_I5914_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5914_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7];
	end
assign N10876 = x_reg_L0_21__retimed_I5914_QOUT;
reg x_reg_L0_21__retimed_I5912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5912_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4];
	end
assign N10869 = x_reg_L0_21__retimed_I5912_QOUT;
reg x_reg_L0_21__retimed_I5911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5911_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4];
	end
assign N10867 = x_reg_L0_21__retimed_I5911_QOUT;
reg x_reg_L0_21__retimed_I5909_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5909_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2];
	end
assign N10860 = x_reg_L0_21__retimed_I5909_QOUT;
reg x_reg_L0_21__retimed_I5908_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5908_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2];
	end
assign N10858 = x_reg_L0_21__retimed_I5908_QOUT;
reg x_reg_L0_21__retimed_I5902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5902_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1];
	end
assign N10841 = x_reg_L0_21__retimed_I5902_QOUT;
reg x_reg_L0_21__retimed_I5901_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5901_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1];
	end
assign N10839 = x_reg_L0_21__retimed_I5901_QOUT;
reg x_reg_L0_21__retimed_I5899_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5899_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6];
	end
assign N10832 = x_reg_L0_21__retimed_I5899_QOUT;
reg x_reg_L0_21__retimed_I5898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5898_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6];
	end
assign N10830 = x_reg_L0_21__retimed_I5898_QOUT;
reg x_reg_L0_21__retimed_I5896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5896_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5];
	end
assign N10823 = x_reg_L0_21__retimed_I5896_QOUT;
reg x_reg_L0_21__retimed_I5895_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5895_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5];
	end
assign N10821 = x_reg_L0_21__retimed_I5895_QOUT;
reg x_reg_L0_21__retimed_I5893_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5893_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0];
	end
assign N10814 = x_reg_L0_21__retimed_I5893_QOUT;
reg x_reg_L0_21__retimed_I5892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5892_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0];
	end
assign N10812 = x_reg_L0_21__retimed_I5892_QOUT;
reg x_reg_L0_21__retimed_I5888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5888_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8];
	end
assign N10800 = x_reg_L0_21__retimed_I5888_QOUT;
reg x_reg_L0_21__retimed_I5887_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5887_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8];
	end
assign N10798 = x_reg_L0_21__retimed_I5887_QOUT;
reg x_reg_L0_21__retimed_I5885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5885_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9];
	end
assign N10792 = x_reg_L0_21__retimed_I5885_QOUT;
reg x_reg_L0_21__retimed_I5884_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5884_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9];
	end
assign N10790 = x_reg_L0_21__retimed_I5884_QOUT;
reg x_reg_L0_21__retimed_I5869_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5869_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27;
	end
assign N10753 = x_reg_L0_21__retimed_I5869_QOUT;
reg x_reg_L0_21__retimed_I5868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5868_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28;
	end
assign N10751 = x_reg_L0_21__retimed_I5868_QOUT;
reg x_reg_L1_21__retimed_I5842_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5842_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44;
	end
assign N10645 = x_reg_L1_21__retimed_I5842_QOUT;
reg x_reg_L1_21__retimed_I5840_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5840_QOUT <= N9758;
	end
assign N10619 = x_reg_L1_21__retimed_I5840_QOUT;
reg x_reg_L1_21__retimed_I5838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5838_QOUT <= N9732;
	end
assign N10593 = x_reg_L1_21__retimed_I5838_QOUT;
reg x_reg_L1_21__retimed_I5836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5836_QOUT <= N9706;
	end
assign N10567 = x_reg_L1_21__retimed_I5836_QOUT;
reg x_reg_L1_21__retimed_I5789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5789_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45];
	end
assign N10428 = x_reg_L1_21__retimed_I5789_QOUT;
reg x_reg_L1_21__retimed_I5786_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5786_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21];
	end
assign N10422 = x_reg_L1_21__retimed_I5786_QOUT;
reg x_reg_L1_20__retimed_I5785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5785_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44];
	end
assign N10419 = x_reg_L1_20__retimed_I5785_QOUT;
reg x_reg_L1_20__retimed_I5782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5782_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20];
	end
assign N10413 = x_reg_L1_20__retimed_I5782_QOUT;
reg x_reg_L1_19__retimed_I5781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5781_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43];
	end
assign N10410 = x_reg_L1_19__retimed_I5781_QOUT;
reg x_reg_L1_19__retimed_I5778_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5778_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19];
	end
assign N10404 = x_reg_L1_19__retimed_I5778_QOUT;
reg x_reg_L1_18__retimed_I5777_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5777_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42];
	end
assign N10401 = x_reg_L1_18__retimed_I5777_QOUT;
reg x_reg_L1_18__retimed_I5774_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5774_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18];
	end
assign N10395 = x_reg_L1_18__retimed_I5774_QOUT;
reg x_reg_L1_17__retimed_I5773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5773_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41];
	end
assign N10392 = x_reg_L1_17__retimed_I5773_QOUT;
reg x_reg_L1_17__retimed_I5770_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5770_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17];
	end
assign N10386 = x_reg_L1_17__retimed_I5770_QOUT;
reg x_reg_L1_16__retimed_I5769_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5769_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40];
	end
assign N10383 = x_reg_L1_16__retimed_I5769_QOUT;
reg x_reg_L1_16__retimed_I5766_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5766_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16];
	end
assign N10377 = x_reg_L1_16__retimed_I5766_QOUT;
reg x_reg_L1_15__retimed_I5765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5765_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39];
	end
assign N10374 = x_reg_L1_15__retimed_I5765_QOUT;
reg x_reg_L1_15__retimed_I5762_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5762_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15];
	end
assign N10368 = x_reg_L1_15__retimed_I5762_QOUT;
reg x_reg_L1_14__retimed_I5761_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5761_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38];
	end
assign N10365 = x_reg_L1_14__retimed_I5761_QOUT;
reg x_reg_L1_14__retimed_I5758_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5758_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N10359 = x_reg_L1_14__retimed_I5758_QOUT;
reg x_reg_L1_13__retimed_I5757_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5757_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37];
	end
assign N10356 = x_reg_L1_13__retimed_I5757_QOUT;
reg x_reg_L1_13__retimed_I5754_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5754_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N10350 = x_reg_L1_13__retimed_I5754_QOUT;
reg x_reg_L1_12__retimed_I5753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5753_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36];
	end
assign N10347 = x_reg_L1_12__retimed_I5753_QOUT;
reg x_reg_L1_12__retimed_I5750_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5750_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N10341 = x_reg_L1_12__retimed_I5750_QOUT;
reg x_reg_L1_11__retimed_I5749_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5749_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35];
	end
assign N10338 = x_reg_L1_11__retimed_I5749_QOUT;
reg x_reg_L1_11__retimed_I5746_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5746_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N10332 = x_reg_L1_11__retimed_I5746_QOUT;
reg x_reg_L1_10__retimed_I5745_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5745_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34];
	end
assign N10329 = x_reg_L1_10__retimed_I5745_QOUT;
reg x_reg_L1_10__retimed_I5742_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5742_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N10323 = x_reg_L1_10__retimed_I5742_QOUT;
reg x_reg_L1_9__retimed_I5741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5741_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33];
	end
assign N10320 = x_reg_L1_9__retimed_I5741_QOUT;
reg x_reg_L1_9__retimed_I5738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5738_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N10314 = x_reg_L1_9__retimed_I5738_QOUT;
reg x_reg_L1_8__retimed_I5737_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5737_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32];
	end
assign N10311 = x_reg_L1_8__retimed_I5737_QOUT;
reg x_reg_L1_8__retimed_I5734_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5734_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N10305 = x_reg_L1_8__retimed_I5734_QOUT;
reg x_reg_L1_7__retimed_I5733_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5733_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31];
	end
assign N10302 = x_reg_L1_7__retimed_I5733_QOUT;
reg x_reg_L1_7__retimed_I5730_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5730_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N10296 = x_reg_L1_7__retimed_I5730_QOUT;
reg x_reg_L1_6__retimed_I5729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5729_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30];
	end
assign N10293 = x_reg_L1_6__retimed_I5729_QOUT;
reg x_reg_L1_6__retimed_I5726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5726_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N10287 = x_reg_L1_6__retimed_I5726_QOUT;
reg x_reg_L1_5__retimed_I5725_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5725_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29];
	end
assign N10284 = x_reg_L1_5__retimed_I5725_QOUT;
reg x_reg_L1_5__retimed_I5722_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5722_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N10278 = x_reg_L1_5__retimed_I5722_QOUT;
reg x_reg_L1_4__retimed_I5721_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5721_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28];
	end
assign N10275 = x_reg_L1_4__retimed_I5721_QOUT;
reg x_reg_L1_4__retimed_I5718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5718_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N10269 = x_reg_L1_4__retimed_I5718_QOUT;
reg x_reg_L1_3__retimed_I5717_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5717_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27];
	end
assign N10266 = x_reg_L1_3__retimed_I5717_QOUT;
reg x_reg_L1_3__retimed_I5714_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5714_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N10260 = x_reg_L1_3__retimed_I5714_QOUT;
reg x_reg_L1_2__retimed_I5713_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5713_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26];
	end
assign N10257 = x_reg_L1_2__retimed_I5713_QOUT;
reg x_reg_L1_2__retimed_I5710_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5710_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N10251 = x_reg_L1_2__retimed_I5710_QOUT;
reg x_reg_L1_1__retimed_I5709_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5709_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25];
	end
assign N10248 = x_reg_L1_1__retimed_I5709_QOUT;
reg x_reg_L1_1__retimed_I5706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5706_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N10242 = x_reg_L1_1__retimed_I5706_QOUT;
reg x_reg_L1_0__retimed_I5705_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5705_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24];
	end
assign N10239 = x_reg_L1_0__retimed_I5705_QOUT;
reg x_reg_L1_0__retimed_I5702_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5702_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N10233 = x_reg_L1_0__retimed_I5702_QOUT;
reg x_reg_L1_21__retimed_I5701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5701_QOUT <= N9257;
	end
assign N10230 = x_reg_L1_21__retimed_I5701_QOUT;
reg x_reg_L1_20__retimed_I5699_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5699_QOUT <= N9252;
	end
assign N10225 = x_reg_L1_20__retimed_I5699_QOUT;
reg x_reg_L1_19__retimed_I5697_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5697_QOUT <= N9247;
	end
assign N10220 = x_reg_L1_19__retimed_I5697_QOUT;
reg x_reg_L1_18__retimed_I5695_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5695_QOUT <= N9242;
	end
assign N10215 = x_reg_L1_18__retimed_I5695_QOUT;
reg x_reg_L1_17__retimed_I5693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5693_QOUT <= N9237;
	end
assign N10210 = x_reg_L1_17__retimed_I5693_QOUT;
reg x_reg_L1_16__retimed_I5691_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5691_QOUT <= N9232;
	end
assign N10205 = x_reg_L1_16__retimed_I5691_QOUT;
reg x_reg_L1_15__retimed_I5689_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5689_QOUT <= N9227;
	end
assign N10200 = x_reg_L1_15__retimed_I5689_QOUT;
reg x_reg_L1_14__retimed_I5687_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5687_QOUT <= N9222;
	end
assign N10195 = x_reg_L1_14__retimed_I5687_QOUT;
reg x_reg_L1_13__retimed_I5685_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5685_QOUT <= N9217;
	end
assign N10190 = x_reg_L1_13__retimed_I5685_QOUT;
reg x_reg_L1_12__retimed_I5683_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5683_QOUT <= N9212;
	end
assign N10185 = x_reg_L1_12__retimed_I5683_QOUT;
reg x_reg_L1_11__retimed_I5681_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5681_QOUT <= N9207;
	end
assign N10180 = x_reg_L1_11__retimed_I5681_QOUT;
reg x_reg_L1_10__retimed_I5679_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5679_QOUT <= N9202;
	end
assign N10175 = x_reg_L1_10__retimed_I5679_QOUT;
reg x_reg_L1_9__retimed_I5677_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5677_QOUT <= N9197;
	end
assign N10170 = x_reg_L1_9__retimed_I5677_QOUT;
reg x_reg_L1_8__retimed_I5675_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5675_QOUT <= N9192;
	end
assign N10165 = x_reg_L1_8__retimed_I5675_QOUT;
reg x_reg_L1_7__retimed_I5673_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5673_QOUT <= N9187;
	end
assign N10160 = x_reg_L1_7__retimed_I5673_QOUT;
reg x_reg_L1_6__retimed_I5671_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5671_QOUT <= N9182;
	end
assign N10155 = x_reg_L1_6__retimed_I5671_QOUT;
reg x_reg_L1_5__retimed_I5669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5669_QOUT <= N9177;
	end
assign N10150 = x_reg_L1_5__retimed_I5669_QOUT;
reg x_reg_L1_4__retimed_I5667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5667_QOUT <= N9172;
	end
assign N10145 = x_reg_L1_4__retimed_I5667_QOUT;
reg x_reg_L1_3__retimed_I5665_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5665_QOUT <= N9167;
	end
assign N10140 = x_reg_L1_3__retimed_I5665_QOUT;
reg x_reg_L1_2__retimed_I5663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5663_QOUT <= N9162;
	end
assign N10135 = x_reg_L1_2__retimed_I5663_QOUT;
reg x_reg_L1_1__retimed_I5661_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5661_QOUT <= N9157;
	end
assign N10130 = x_reg_L1_1__retimed_I5661_QOUT;
reg x_reg_L1_0__retimed_I5659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5659_QOUT <= N9152;
	end
assign N10125 = x_reg_L1_0__retimed_I5659_QOUT;
reg x_reg_L1_21__retimed_I5654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5654_QOUT <= N9141;
	end
assign N10114 = x_reg_L1_21__retimed_I5654_QOUT;
reg x_reg_L1_20__retimed_I5650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5650_QOUT <= N9132;
	end
assign N10105 = x_reg_L1_20__retimed_I5650_QOUT;
reg x_reg_L1_19__retimed_I5646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5646_QOUT <= N9123;
	end
assign N10096 = x_reg_L1_19__retimed_I5646_QOUT;
reg x_reg_L1_18__retimed_I5642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5642_QOUT <= N9114;
	end
assign N10087 = x_reg_L1_18__retimed_I5642_QOUT;
reg x_reg_L1_17__retimed_I5638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5638_QOUT <= N9105;
	end
assign N10078 = x_reg_L1_17__retimed_I5638_QOUT;
reg x_reg_L1_16__retimed_I5634_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5634_QOUT <= N9096;
	end
assign N10069 = x_reg_L1_16__retimed_I5634_QOUT;
reg x_reg_L1_15__retimed_I5630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5630_QOUT <= N9087;
	end
assign N10060 = x_reg_L1_15__retimed_I5630_QOUT;
reg x_reg_L1_14__retimed_I5626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5626_QOUT <= N9078;
	end
assign N10051 = x_reg_L1_14__retimed_I5626_QOUT;
reg x_reg_L1_13__retimed_I5622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5622_QOUT <= N9069;
	end
assign N10042 = x_reg_L1_13__retimed_I5622_QOUT;
reg x_reg_L1_12__retimed_I5618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5618_QOUT <= N9060;
	end
assign N10033 = x_reg_L1_12__retimed_I5618_QOUT;
reg x_reg_L1_11__retimed_I5614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5614_QOUT <= N9051;
	end
assign N10024 = x_reg_L1_11__retimed_I5614_QOUT;
reg x_reg_L1_10__retimed_I5610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5610_QOUT <= N9042;
	end
assign N10015 = x_reg_L1_10__retimed_I5610_QOUT;
reg x_reg_L1_9__retimed_I5606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5606_QOUT <= N9033;
	end
assign N10006 = x_reg_L1_9__retimed_I5606_QOUT;
reg x_reg_L1_8__retimed_I5602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5602_QOUT <= N9024;
	end
assign N9997 = x_reg_L1_8__retimed_I5602_QOUT;
reg x_reg_L1_7__retimed_I5598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5598_QOUT <= N9015;
	end
assign N9988 = x_reg_L1_7__retimed_I5598_QOUT;
reg x_reg_L1_6__retimed_I5594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5594_QOUT <= N9006;
	end
assign N9979 = x_reg_L1_6__retimed_I5594_QOUT;
reg x_reg_L1_5__retimed_I5590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5590_QOUT <= N8997;
	end
assign N9970 = x_reg_L1_5__retimed_I5590_QOUT;
reg x_reg_L1_4__retimed_I5586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5586_QOUT <= N8988;
	end
assign N9961 = x_reg_L1_4__retimed_I5586_QOUT;
reg x_reg_L1_3__retimed_I5582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5582_QOUT <= N8979;
	end
assign N9952 = x_reg_L1_3__retimed_I5582_QOUT;
reg x_reg_L1_2__retimed_I5578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5578_QOUT <= N8970;
	end
assign N9943 = x_reg_L1_2__retimed_I5578_QOUT;
reg x_reg_L1_1__retimed_I5574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5574_QOUT <= N8961;
	end
assign N9934 = x_reg_L1_1__retimed_I5574_QOUT;
reg x_reg_L1_0__retimed_I5573_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5573_QOUT <= N8958;
	end
assign N9931 = x_reg_L1_0__retimed_I5573_QOUT;
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6872 (.Y(N13249), .A(N9931));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6873 (.Y(N13250), .A(N13249));
reg x_reg_L1_0__retimed_I5570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5570_QOUT <= N8952;
	end
assign N9925 = x_reg_L1_0__retimed_I5570_QOUT;
reg x_reg_L0_21__retimed_I5520_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5520_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26;
	end
assign N9758 = x_reg_L0_21__retimed_I5520_QOUT;
reg x_reg_L0_21__retimed_I5518_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5518_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144;
	end
assign N9732 = x_reg_L0_21__retimed_I5518_QOUT;
reg x_reg_L0_21__retimed_I5516_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5516_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225;
	end
assign N9706 = x_reg_L0_21__retimed_I5516_QOUT;
reg x_reg_L1_22__retimed_I5514_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5514_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053;
	end
assign N9680 = x_reg_L1_22__retimed_I5514_QOUT;
reg x_reg_L1_22__retimed_I5513_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5513_QOUT <= N8945;
	end
assign N9678 = x_reg_L1_22__retimed_I5513_QOUT;
reg x_reg_L1_23__retimed_I5511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5511_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004;
	end
assign N9673 = x_reg_L1_23__retimed_I5511_QOUT;
reg x_reg_L1_23__retimed_I5510_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5510_QOUT <= N8938;
	end
assign N9671 = x_reg_L1_23__retimed_I5510_QOUT;
reg x_reg_L1_24__retimed_I5508_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__retimed_I5508_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1];
	end
assign N9666 = x_reg_L1_24__retimed_I5508_QOUT;
reg x_reg_L1_25__retimed_I5505_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__retimed_I5505_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2];
	end
assign N9659 = x_reg_L1_25__retimed_I5505_QOUT;
reg x_reg_L1_26__retimed_I5502_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__retimed_I5502_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3];
	end
assign N9652 = x_reg_L1_26__retimed_I5502_QOUT;
reg x_reg_L1_27__retimed_I5499_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__retimed_I5499_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4];
	end
assign N9645 = x_reg_L1_27__retimed_I5499_QOUT;
reg x_reg_L1_28__retimed_I5496_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__retimed_I5496_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5];
	end
assign N9638 = x_reg_L1_28__retimed_I5496_QOUT;
reg x_reg_L1_29__retimed_I5494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I5494_QOUT <= N8900;
	end
assign N9633 = x_reg_L1_29__retimed_I5494_QOUT;
reg x_reg_L1_29__retimed_I5493_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I5493_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6];
	end
assign N9631 = x_reg_L1_29__retimed_I5493_QOUT;
reg x_reg_L1_30__retimed_I5490_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__retimed_I5490_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7];
	end
assign N9624 = x_reg_L1_30__retimed_I5490_QOUT;
reg x_reg_L0_21__retimed_I5330_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5330_QOUT <= a_man[21];
	end
assign N9257 = x_reg_L0_21__retimed_I5330_QOUT;
reg x_reg_L0_20__retimed_I5328_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5328_QOUT <= a_man[20];
	end
assign N9252 = x_reg_L0_20__retimed_I5328_QOUT;
reg x_reg_L0_19__retimed_I5326_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5326_QOUT <= a_man[19];
	end
assign N9247 = x_reg_L0_19__retimed_I5326_QOUT;
reg x_reg_L0_18__retimed_I5324_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5324_QOUT <= a_man[18];
	end
assign N9242 = x_reg_L0_18__retimed_I5324_QOUT;
reg x_reg_L0_17__retimed_I5322_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5322_QOUT <= a_man[17];
	end
assign N9237 = x_reg_L0_17__retimed_I5322_QOUT;
reg x_reg_L0_16__retimed_I5320_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5320_QOUT <= a_man[16];
	end
assign N9232 = x_reg_L0_16__retimed_I5320_QOUT;
reg x_reg_L0_15__retimed_I5318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5318_QOUT <= a_man[15];
	end
assign N9227 = x_reg_L0_15__retimed_I5318_QOUT;
reg x_reg_L0_14__retimed_I5316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5316_QOUT <= a_man[14];
	end
assign N9222 = x_reg_L0_14__retimed_I5316_QOUT;
reg x_reg_L0_13__retimed_I5314_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5314_QOUT <= a_man[13];
	end
assign N9217 = x_reg_L0_13__retimed_I5314_QOUT;
reg x_reg_L0_12__retimed_I5312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5312_QOUT <= a_man[12];
	end
assign N9212 = x_reg_L0_12__retimed_I5312_QOUT;
reg x_reg_L0_11__retimed_I5310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5310_QOUT <= a_man[11];
	end
assign N9207 = x_reg_L0_11__retimed_I5310_QOUT;
reg x_reg_L0_10__retimed_I5308_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5308_QOUT <= a_man[10];
	end
assign N9202 = x_reg_L0_10__retimed_I5308_QOUT;
reg x_reg_L0_9__retimed_I5306_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5306_QOUT <= a_man[9];
	end
assign N9197 = x_reg_L0_9__retimed_I5306_QOUT;
reg x_reg_L0_8__retimed_I5304_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5304_QOUT <= a_man[8];
	end
assign N9192 = x_reg_L0_8__retimed_I5304_QOUT;
reg x_reg_L0_7__retimed_I5302_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5302_QOUT <= a_man[7];
	end
assign N9187 = x_reg_L0_7__retimed_I5302_QOUT;
reg x_reg_L0_6__retimed_I5300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5300_QOUT <= a_man[6];
	end
assign N9182 = x_reg_L0_6__retimed_I5300_QOUT;
reg x_reg_L0_5__retimed_I5298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5298_QOUT <= a_man[5];
	end
assign N9177 = x_reg_L0_5__retimed_I5298_QOUT;
reg x_reg_L0_4__retimed_I5296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5296_QOUT <= a_man[4];
	end
assign N9172 = x_reg_L0_4__retimed_I5296_QOUT;
reg x_reg_L0_3__retimed_I5294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5294_QOUT <= a_man[3];
	end
assign N9167 = x_reg_L0_3__retimed_I5294_QOUT;
reg x_reg_L0_2__retimed_I5292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5292_QOUT <= a_man[2];
	end
assign N9162 = x_reg_L0_2__retimed_I5292_QOUT;
reg x_reg_L0_1__retimed_I5290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5290_QOUT <= a_man[1];
	end
assign N9157 = x_reg_L0_1__retimed_I5290_QOUT;
reg x_reg_L0_0__retimed_I5288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5288_QOUT <= a_man[0];
	end
assign N9152 = x_reg_L0_0__retimed_I5288_QOUT;
reg x_reg_L0_21__retimed_I5283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5283_QOUT <= b_man[21];
	end
assign N9141 = x_reg_L0_21__retimed_I5283_QOUT;
reg x_reg_L0_20__retimed_I5279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5279_QOUT <= b_man[20];
	end
assign N9132 = x_reg_L0_20__retimed_I5279_QOUT;
reg x_reg_L0_19__retimed_I5275_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5275_QOUT <= b_man[19];
	end
assign N9123 = x_reg_L0_19__retimed_I5275_QOUT;
reg x_reg_L0_18__retimed_I5271_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5271_QOUT <= b_man[18];
	end
assign N9114 = x_reg_L0_18__retimed_I5271_QOUT;
reg x_reg_L0_17__retimed_I5267_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5267_QOUT <= b_man[17];
	end
assign N9105 = x_reg_L0_17__retimed_I5267_QOUT;
reg x_reg_L0_16__retimed_I5263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5263_QOUT <= b_man[16];
	end
assign N9096 = x_reg_L0_16__retimed_I5263_QOUT;
reg x_reg_L0_15__retimed_I5259_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5259_QOUT <= b_man[15];
	end
assign N9087 = x_reg_L0_15__retimed_I5259_QOUT;
reg x_reg_L0_14__retimed_I5255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5255_QOUT <= b_man[14];
	end
assign N9078 = x_reg_L0_14__retimed_I5255_QOUT;
reg x_reg_L0_13__retimed_I5251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5251_QOUT <= b_man[13];
	end
assign N9069 = x_reg_L0_13__retimed_I5251_QOUT;
reg x_reg_L0_12__retimed_I5247_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5247_QOUT <= b_man[12];
	end
assign N9060 = x_reg_L0_12__retimed_I5247_QOUT;
reg x_reg_L0_11__retimed_I5243_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5243_QOUT <= b_man[11];
	end
assign N9051 = x_reg_L0_11__retimed_I5243_QOUT;
reg x_reg_L0_10__retimed_I5239_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5239_QOUT <= b_man[10];
	end
assign N9042 = x_reg_L0_10__retimed_I5239_QOUT;
reg x_reg_L0_9__retimed_I5235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5235_QOUT <= b_man[9];
	end
assign N9033 = x_reg_L0_9__retimed_I5235_QOUT;
reg x_reg_L0_8__retimed_I5231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5231_QOUT <= b_man[8];
	end
assign N9024 = x_reg_L0_8__retimed_I5231_QOUT;
reg x_reg_L0_7__retimed_I5227_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5227_QOUT <= b_man[7];
	end
assign N9015 = x_reg_L0_7__retimed_I5227_QOUT;
reg x_reg_L0_6__retimed_I5223_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5223_QOUT <= b_man[6];
	end
assign N9006 = x_reg_L0_6__retimed_I5223_QOUT;
reg x_reg_L0_5__retimed_I5219_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5219_QOUT <= b_man[5];
	end
assign N8997 = x_reg_L0_5__retimed_I5219_QOUT;
reg x_reg_L0_4__retimed_I5215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5215_QOUT <= b_man[4];
	end
assign N8988 = x_reg_L0_4__retimed_I5215_QOUT;
reg x_reg_L0_3__retimed_I5211_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5211_QOUT <= b_man[3];
	end
assign N8979 = x_reg_L0_3__retimed_I5211_QOUT;
reg x_reg_L0_2__retimed_I5207_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5207_QOUT <= b_man[2];
	end
assign N8970 = x_reg_L0_2__retimed_I5207_QOUT;
reg x_reg_L0_1__retimed_I5203_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5203_QOUT <= b_man[1];
	end
assign N8961 = x_reg_L0_1__retimed_I5203_QOUT;
reg x_reg_L0_0__retimed_I5202_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5202_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47;
	end
assign N8958 = x_reg_L0_0__retimed_I5202_QOUT;
reg x_reg_L0_0__retimed_I5199_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5199_QOUT <= b_man[0];
	end
assign N8952 = x_reg_L0_0__retimed_I5199_QOUT;
reg x_reg_L0_22__retimed_I5196_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5196_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055;
	end
assign N8945 = x_reg_L0_22__retimed_I5196_QOUT;
reg x_reg_L0_23__retimed_I5193_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I5193_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025;
	end
assign N8938 = x_reg_L0_23__retimed_I5193_QOUT;
reg x_reg_L0_29__retimed_I5177_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__retimed_I5177_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008;
	end
assign N8900 = x_reg_L0_29__retimed_I5177_QOUT;
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007), .A(a_exp[0]), .B(a_exp[1]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I2 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I3 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434), .A(a_exp[7]), .B(a_exp[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2009));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I4 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2007), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8434));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I5 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2043));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I7 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I8 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I9 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I10 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I11 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2030), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2049), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2038), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2058));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I12 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I13 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I14 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2041), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2052), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2062));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I15 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I16 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896), .A(b_exp[0]), .B(b_exp[1]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I17 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I18 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426), .A(b_exp[7]), .B(b_exp[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1898));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I19 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1896), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8426));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I20 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I21 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1932));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I22 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919), .A(b_man[10]), .B(b_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I23 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938), .A(b_man[6]), .B(b_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I24 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927), .A(b_man[8]), .B(b_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I25 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947), .A(b_man[4]), .B(b_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I26 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1919), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1938), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1927), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1947));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I27 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I28 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I29 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1936), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1930), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1941), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1951));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I30 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I31 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I32 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I33 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I34 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I35 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1981), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1988), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1985), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N1976));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I36 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__19));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I37 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I38 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092), .A(b_exp[0]), .B(b_exp[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I39 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099), .A(b_exp[5]), .B(b_exp[4]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I40 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096), .A(b_exp[7]), .B(b_exp[6]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I41 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087), .A(b_exp[3]), .B(b_exp[2]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I42 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2092), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2099), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2096), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2087));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I43 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__12));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I44 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I45 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N441), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N440));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I46 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6225), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I47 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0]), .A(b_exp[0]), .B(a_exp[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I48 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[0]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I49 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .A(b_man[22]), .B(b_man[21]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I50 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I51 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .A(a_man[22]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I52 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .A(a_man[20]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I53 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I54 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .A(a_man[21]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I55 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I56 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I57 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011), .A(b_man[22]), .B(b_man[21]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I58 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I59 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2466));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I60 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3183), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2327));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I61 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .A(b_man[20]), .B(b_man[19]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I62 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007), .A(b_man[21]), .B(b_man[19]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I63 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3007), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I64 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552), .A(b_man[21]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I65 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I66 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2183));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I67 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .A(a_man[18]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I68 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I69 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .A(a_man[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I70 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I71 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I72 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2675));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I73 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3726), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3039), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I74 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I75 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2964), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3380), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2703));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I76 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2998), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3110), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2851));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I77 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3166), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I78 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I79 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I80 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I81 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3640), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I82 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .A(a_man[16]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I83 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I84 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .A(a_man[17]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I85 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I86 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I87 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2884));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I88 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2313), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3241), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I89 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I90 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3568), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3580), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3296));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I91 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3305), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2603), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3712));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I92 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2755), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2381), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2391));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I93 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I94 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169), .A(b_man[19]), .B(b_man[17]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I95 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .A(b_man[18]), .B(b_man[17]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I96 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2169), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I97 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407), .A(b_man[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I98 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I99 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I101 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2955), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I102 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2455), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2592), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3371));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I103 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I104 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2250));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I105 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2249), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2632), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3181));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I107 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3367));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .A(b_man[16]), .B(b_man[15]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973), .A(b_man[17]), .B(b_man[15]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I110 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2973), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268), .A(b_man[17]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2309));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .A(a_man[14]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I115 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I116 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .A(a_man[15]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I117 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I118 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I119 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3095));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2526), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3438), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I122 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3686), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2177), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2534));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I126 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I127 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I128 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I129 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I131 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2809), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2662), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2522));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I132 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2275), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3287), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3086));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I133 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2241), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3160), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3711), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3030), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I135 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3503), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3372), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2409));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I136 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3029), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3230), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3437));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I137 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2170), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I140 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I141 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2301), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I142 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3434), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3344), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3569));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I143 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3143), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2935), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2729));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I144 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2515), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2873), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2146));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I145 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I146 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3333), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3564));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I147 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .A(a_man[12]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I149 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .A(a_man[13]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I152 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3297));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2740), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3634), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I154 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I155 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2197), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2374), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3650));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I156 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I157 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2447), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I158 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I160 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I162 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I164 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .A(a_man[10]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I165 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I166 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .A(a_man[11]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I169 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3496));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I170 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2949), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2232), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I171 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I172 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3433), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2587), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3431));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I173 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2295), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2163), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2462));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I175 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I177 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124), .A(b_man[15]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I178 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I179 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .A(b_man[14]), .B(b_man[13]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751), .A(b_man[15]), .B(b_man[13]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I182 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3751), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I183 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I184 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3631), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3499), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3058));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I185 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2234));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I186 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3092), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2369), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I187 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3229), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2516), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I188 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2590), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2734), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2874));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I189 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3457), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2190));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I190 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3398), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3704), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3203));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I191 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I192 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2376));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I193 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3540), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3543), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3279));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I194 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2576), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2792), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2681));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I195 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I196 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3366), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2654), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I197 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .A(b_man[12]), .B(b_man[11]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I198 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942), .A(b_man[13]), .B(b_man[11]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I199 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2942), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I200 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981), .A(b_man[13]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I201 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I202 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2451));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I203 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I204 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3292), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I205 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I206 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3156), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I207 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I209 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2945), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2803), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2658));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I210 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3201), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2256), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2790));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I211 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3060), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3023), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2906));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I212 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2427), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3000), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3021));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I213 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I214 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2161));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I215 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I216 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3562), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I217 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I218 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3427), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I219 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3222), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3087), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3719));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I220 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I221 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2296), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I222 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I223 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2443), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I224 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3091), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3700));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I225 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2880), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3515), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3575));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I226 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3116), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3320), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2970));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I227 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2846), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2697), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3532));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I228 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I229 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I230 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I231 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I232 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I233 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I234 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I235 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I236 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I238 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3286), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3150), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3419));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720), .A(b_man[11]), .B(b_man[9]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .A(b_man[10]), .B(b_man[9]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3720), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I242 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827), .A(b_man[11]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I244 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I246 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3224), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I247 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I248 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3359), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I249 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2732), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2868), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3018));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I250 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3293), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2230), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2823));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I251 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2728), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3626), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I252 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2583), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3492), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I253 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2865), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2157), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I254 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2363), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2228), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2508));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I255 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .A(a_man[8]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I257 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .A(a_man[9]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I258 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I259 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I260 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3699));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I261 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3153), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2440), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I262 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I263 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3066), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2801), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3469));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2518));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I266 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3692), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2843), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2556));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I267 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2308), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3576));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I268 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2551), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2762), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2514));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I270 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2360));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3527));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I273 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2797), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I275 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2650), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I276 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2936), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I278 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2436), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2290), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2577));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I280 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2511), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2364), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I283 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2160), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3629), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3136));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I284 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2496), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2705), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3612));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I285 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .A(a_man[6]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .A(a_man[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I288 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I289 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I290 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2289));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I291 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3356), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2647), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I292 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I293 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2179), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3015), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2165));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I294 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I295 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3081), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .A(b_man[8]), .B(b_man[7]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911), .A(b_man[9]), .B(b_man[7]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678), .A(b_man[9]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I300 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I301 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2586));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I302 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2720), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2487));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I303 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3550), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3358));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I304 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3491), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2944), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2172));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I305 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3377), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2611), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3318));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I306 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I307 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I308 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3693), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I309 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I310 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3559), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I311 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I312 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2222), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I313 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3350), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3216), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3486));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3421), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I317 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3289), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I318 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I319 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I320 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3084), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2937), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2799));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I321 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3122), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3666), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2867));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I322 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2582), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3753), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3149));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I323 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3235), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2736), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2283));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2571));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I326 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I327 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2356), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I328 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3520), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3622), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3326));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I329 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .A(a_man[4]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I330 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I331 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .A(a_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I332 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I333 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I334 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2500));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I335 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3555), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2858), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I336 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I337 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2923), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3214), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2743));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I338 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .A(b_man[6]), .B(b_man[5]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I339 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691), .A(b_man[7]), .B(b_man[5]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I340 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3691), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531), .A(b_man[7]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2653));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I345 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2860), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2723), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I349 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3010), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I350 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2503), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2359), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2642));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I351 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3017), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3744), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3177));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I353 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2149), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I354 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3624), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2284), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I358 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3412), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3283), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3551));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I360 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I362 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I366 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I367 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2863), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3013), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3147));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I368 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2439), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3354), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I369 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2580), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3487), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I370 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3698), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3441), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2225));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I371 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2589), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3155), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3435));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I372 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2315), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2887), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3653));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I373 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3406), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2557), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2202));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I374 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2677), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3243), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2302));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I375 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2770), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2343), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2596));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I376 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3009), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3210), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3097));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I377 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I378 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I379 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3281), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I380 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3144), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I382 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I384 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I385 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3211), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I388 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I389 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I390 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3001), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2853), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3135));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I391 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2649), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3414), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2617));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I392 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2927), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2791), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2236));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I393 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3728), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2405), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3464));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I394 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2855), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3606), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2320));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I396 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2787));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I397 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3413), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3733));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I398 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2570), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3477), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I399 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2428), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3345), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I400 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I401 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I406 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I407 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I409 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3479), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3347), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3615));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I411 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I412 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I413 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I414 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881), .A(b_man[5]), .B(b_man[3]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .A(b_man[4]), .B(b_man[3]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2881), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377), .A(b_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I420 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I421 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I422 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3213), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3078), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2933));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I423 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2929), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2218), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2794), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3690), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I425 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3075), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2349), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I426 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2429), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2714));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I427 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2477), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2387));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I428 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2216), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3687), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3614));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I429 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3636), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2908));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2645), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3554), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I431 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2506), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3416), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I432 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2288), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2154), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2660));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I433 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2351), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2564), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2889));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I434 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .A(a_man[2]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I435 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I436 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .A(a_man[3]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I437 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I438 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I439 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2711));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I440 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2147), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3071), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I441 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I442 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3164), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3410), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3572));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I443 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I446 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3274), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I449 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I450 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I451 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3067), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2921), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3204));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3003), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I454 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I455 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2857), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I456 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I457 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3140), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I458 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2639), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2498), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2786));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I459 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3104), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3644), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3715));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I460 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2210), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2686), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3192));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I461 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2442), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2861), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2344));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I462 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3583), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2804), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3300));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I463 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3382), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3186), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3393));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I464 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I465 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I466 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2726));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I467 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2635), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3541), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I468 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2497), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3404), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I469 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I470 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2783), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I471 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2278), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3754), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2421));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I472 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3396), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2987), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3736));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I473 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I474 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2718), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014), .A(b_man[2]), .B(b_man[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6874 (.Y(N13251), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6875 (.Y(N13252), .A(N13251));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662), .A(b_man[3]), .B(b_man[1]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I477 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3662), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3014));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I478 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237), .A(b_man[3]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796), .A0(N13252), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I480 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2796));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2347), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .A(a_man[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I483 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I485 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3611), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3079));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I486 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I487 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2575), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I488 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2812), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2931), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2221));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I489 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2353), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3057), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3494));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I490 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I491 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2144), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I492 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I493 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3619), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I494 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I495 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2280), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I496 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3409), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3278), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3544));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I498 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3483), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357), .B(N13252), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I501 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3142), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2572), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3008));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I502 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2510), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3083), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3239));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I503 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2245), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3734), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3309));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I504 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3273), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2416), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3474));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I505 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3498), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3074), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2502));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I506 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3042), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3098), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2636));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I507 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I508 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I509 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2321), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2597), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3455));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I510 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I511 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I512 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I513 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I515 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I516 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I517 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I518 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I519 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3267), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3534));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I520 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I522 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I524 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3207), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I525 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I527 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I528 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2849), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3130));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I529 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3339), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2272), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2953));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I530 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2925), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I533 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2789), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I534 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I535 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3068), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I536 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2568), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2425), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2710));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I537 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2640), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I539 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3271), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I540 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I541 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2282), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2919), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2845));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I542 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2840), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2693), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3220));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I543 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I544 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2271), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I545 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2847), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3747), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I546 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2565), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3470), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2422), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3340), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I548 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2706), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3607), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I549 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2211), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3682), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2341));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I550 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2628), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2488), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2682));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I551 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2159), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2722), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3223));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I552 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2833), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2540), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3200));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I553 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2622), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3673));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I554 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2950), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2291), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3696));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I555 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I556 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3679), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2991), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I557 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3337), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3565), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2976));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I558 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .A(b_man[0]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I559 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361), .A(b_man[1]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I561 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I562 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2859));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I563 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2695), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2454));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I565 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2346), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I567 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2214), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I568 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I569 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2489), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I570 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3608), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3475), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3750));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I571 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I573 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3548), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I575 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I576 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3684), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I577 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3070), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3209), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3343));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I578 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3657), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2607), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2999));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I579 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2562), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .A(a_man[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I581 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I582 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3467), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I583 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831), .A(b_man[21]), .B(b_man[22]));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I584 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I585 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2831), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2411));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I586 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3128), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2492));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I587 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2206), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2775), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3628));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I588 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2778), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I590 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2631), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I592 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I593 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2913), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I594 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2414), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2273), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2558));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I595 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3174), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3113), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2727));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I596 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2996), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2484), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3538));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I597 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2959), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3026), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2702));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I598 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2265), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2752), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2186));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I599 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2148), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3472), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3218));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I600 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I601 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I602 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I603 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I604 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3133), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I605 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I606 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2997), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I607 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I608 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3270), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I609 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2781), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2633), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2917));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I610 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I611 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2712), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I612 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I613 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2852), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I614 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2348), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3288), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2493));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I615 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2517), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3088), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2769));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I616 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I617 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3674), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I618 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I619 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3536), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I620 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I621 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2203), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I622 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3332), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3199), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3463));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I623 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3570), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2494));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I624 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I625 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3196), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I626 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I627 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3059), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I628 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2839), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2698), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2227));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I629 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2253), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3315), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2758));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I630 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2361), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2785), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2410));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I631 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2385), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3506), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2657));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I632 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3331), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3590), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2932));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I633 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I634 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I635 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3401), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I636 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I637 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2841), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I638 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I639 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2701), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I640 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I641 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2985), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I642 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2482), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2338), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2623));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I643 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3061), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2432), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2208));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I644 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I645 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2419), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I646 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I647 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2276), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I648 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I649 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2559), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I650 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3677), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3539), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2205));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I651 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2862), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I652 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3610), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I653 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I654 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3752), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I655 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3272), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3749), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3403));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I656 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3006), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3547), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2473));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I657 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I658 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2480), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I659 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I660 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2335), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I661 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3739), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3599), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3556));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I662 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2166), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2731), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3233));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I663 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2630), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2547), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2191));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I664 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2870), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3423), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2424));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I665 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2450), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2433));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I666 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I667 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3395));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I668 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2504), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I669 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2920), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I670 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I671 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3065), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I672 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2561), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2704));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I673 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I674 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I675 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I676 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I677 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I678 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I679 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I680 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I681 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I682 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2198), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3667), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2328));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I683 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3322), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2909), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3535));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I684 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I685 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3742), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I686 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I687 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3601), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I688 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I689 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2266), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I690 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3264), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3526));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I691 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I692 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3336), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I693 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I694 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3202), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I695 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I696 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3466), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I697 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2844), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3125));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I698 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3459), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2402), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2192));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I699 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3261), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2549), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I700 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3123), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2406), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I701 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2907), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2771), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3282));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I702 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2638), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3206), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3689));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I703 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3510), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3031), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3574));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I704 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3198), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3741), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2194));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I705 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2298), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2217), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2145));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I706 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I707 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I708 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2910), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I709 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I710 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2774), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I711 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I712 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3054), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I713 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2408), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2694));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I714 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I715 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2485), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I716 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I717 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2340), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I718 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I719 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2626), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I720 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3745), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3605), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2270));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I721 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2673), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3238), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3262));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I722 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3392), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2691), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I723 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I724 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3327), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I725 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I726 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3193), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I727 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I728 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3458), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I729 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2979), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2834), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3115));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I730 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2974), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3723), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3002));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I731 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3119), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3053), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2554));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I732 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2366), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3490), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I733 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2393), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2965), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2666));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I734 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3681), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3597), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3533));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I735 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I736 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3596));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I737 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2539));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I738 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3016), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3613));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I739 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543), .A(b_man[19]), .B(b_man[20]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I740 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901), .A(b_man[21]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2543));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I741 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2152), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I742 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2207), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I743 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2901), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3468));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I744 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I745 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2330), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I746 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I747 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2200), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I748 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I749 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2474), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I750 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3595), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3460), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3735));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I751 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I752 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3531), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I753 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I754 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3397), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I755 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I756 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3668), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I757 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3194), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3056), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3329));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I758 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2947), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3493), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2708));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I759 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3664), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2525), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2311));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I760 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2848), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2337), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3024));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I761 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2876), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3429), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3146));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I762 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2457), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3319));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I763 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I764 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2199), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2765), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2730));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I765 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3346), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2279), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3604));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I766 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2304), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2939), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3041));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I767 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I768 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I769 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I770 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2763), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I771 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I772 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2616), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I773 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610), .A(b_man[17]), .B(b_man[18]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I774 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971), .A(b_man[19]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2610));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I775 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3415), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I776 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3076), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I777 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I778 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2971), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3671));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I779 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2400), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2261), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2345));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I780 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3593), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2392), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3552), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2756));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I781 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2370), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3255), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2882));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I782 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3127), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2412), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I783 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I784 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3265), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I785 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2776), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2912));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I786 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2438), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2175), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2437));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I787 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I788 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3521), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I789 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I790 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3387), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I791 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3659), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2463), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3407), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2819));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I792 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3184), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3048), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3321));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I793 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2287), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3500));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I794 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I795 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3117), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I796 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I797 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2983), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I798 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I799 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3258), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I800 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2766), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2618), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2903));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I801 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I802 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2696), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I803 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I804 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2555), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I805 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I806 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2837), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I807 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2332), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2201), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2479));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I808 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2856), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3408), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2151));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I809 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2585), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3152), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2173));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I810 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3180), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3378), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2820));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I811 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3400), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2793), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2748));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I812 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I813 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2716), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I814 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3330), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I815 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I816 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3462), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I817 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2984), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3120));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I818 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2619), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3609), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2961));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I819 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I820 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2545), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I821 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I822 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2403), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I823 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I824 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2687), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I825 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2195), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3661), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2322));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I826 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I827 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3737), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I828 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I829 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3598), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I830 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I831 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2263), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I832 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3259), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3524));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I833 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2773), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3328), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3226));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I834 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3069), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3244));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I835 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3037), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3578), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3633));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I836 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2614), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3263), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2456));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I837 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I838 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2396));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I839 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2922), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2751));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I840 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I841 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3323), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I842 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I843 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3187), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I844 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I845 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3453), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I846 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2975), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2829), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3111));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I847 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I848 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2905), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I849 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I850 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2768), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I851 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I852 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3052), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I853 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2548), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2404), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2689));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I854 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3045), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3584), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2397));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I855 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676), .A(b_man[15]), .B(b_man[16]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I856 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043), .A(b_man[17]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2676));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I857 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I858 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2620), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I859 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3043), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2264));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I860 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I861 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2826), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I862 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2890), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2469), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2262));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I863 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2407), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2204), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2688));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I864 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2231), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2800), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3553));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I865 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3436), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2464), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3516));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I866 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I867 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3727), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2529), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3268), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2888));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I868 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I869 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3587), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I870 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I871 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3525), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I872 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I873 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3665), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I874 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3190), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3324));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I875 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3383), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3251), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2238));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I876 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2470), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2982), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3743));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I877 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3465), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2709), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2143));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I878 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3295), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3355), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2980));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I879 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I880 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I881 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2532), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3246), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2940));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I882 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I883 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2759), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I884 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I885 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2612), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I886 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I887 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2895), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I888 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2258), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2537));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I889 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I890 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2326), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I891 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I892 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2196), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I893 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I894 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2471), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I895 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3592), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3456), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3729));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I896 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2745), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3302), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3208));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I897 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3730), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2680), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3670));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I898 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3269), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3212), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2418));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I899 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749), .A(b_man[13]), .B(b_man[14]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I900 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105), .A(b_man[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2749));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I901 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I902 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2832), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I903 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3105), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2472));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I904 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3219), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3501), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3724));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I905 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I906 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3518), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I907 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I908 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3385), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I909 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I910 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3654), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I911 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3046), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3316));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I912 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I913 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3114), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I914 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I915 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2978), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I916 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I917 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3252), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I918 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2760), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2615), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2898));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I919 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3702), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2652), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2372));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I920 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2378), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2951), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2316));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I921 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3126), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3523), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3482));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I922 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I923 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I924 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2187), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2598), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3124), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2960));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I925 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2924), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I926 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3731), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I927 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I928 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2259), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I929 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3386), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3519));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I930 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3448), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2926), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2918));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I931 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I932 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2542), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I933 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I934 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2398), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I935 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I936 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2679), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I937 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2188), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3658), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2317));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I938 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2864), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3618), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3189));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I939 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3363), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2292), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2591));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I940 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3384), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2181), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2667));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I941 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I942 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I943 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3317), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I944 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I945 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3182), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I946 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I947 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3451), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I948 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2969), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2822), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3109));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I949 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I950 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2966), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I951 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I952 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2821), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I953 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817), .A(b_man[11]), .B(b_man[12]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I954 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172), .A(b_man[13]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2817));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I955 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I956 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3047), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I957 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3172), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2683));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I958 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2604), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2465), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2625));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I959 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3335), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3277), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3703));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I960 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2717), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3077), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3560));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I961 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3638), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3158), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3461));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I962 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I963 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I964 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I965 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I966 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3721), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I967 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I968 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3585), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I969 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2254), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2664), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2981), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3032));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I970 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3379), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3245), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3511));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I971 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I972 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2753), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I973 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I974 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2608), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I975 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I976 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2891), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I977 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2390), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2255), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2533));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I978 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2269), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2478), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2627));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I979 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2780), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2567), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2420));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I980 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3020), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2505), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2646));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I981 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I982 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I983 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2319), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I984 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I985 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2467), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I986 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3586), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3725));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I987 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883), .A(b_man[9]), .B(b_man[10]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I988 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236), .A(b_man[11]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2883));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I989 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I990 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3247), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I991 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3236), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2892));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I992 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I993 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3038), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I994 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2312), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2737), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2827), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3094));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I995 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I996 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2180), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I997 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3131), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I998 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2535), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I999 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1000 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1001 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1002 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2182), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2314));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1003 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3579), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3443), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2601));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1004 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3450), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2671), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2325));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1005 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2989), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3051), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3530));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1006 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2213), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2354), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3444));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1007 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1008 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1009 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1010 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3514), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1011 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3381), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2674), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1012 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1013 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3648), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1014 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3175), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3040), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3310));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1015 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2897), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3170));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1016 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3738), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3676), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2355));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1017 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1018 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1019 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2963), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1020 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1021 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2818), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1022 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1023 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3101), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1024 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2602), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2461), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2744));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1025 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3108), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3311), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3685));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1026 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3390), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2541), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2899));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1027 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1028 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952), .A(b_man[7]), .B(b_man[8]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1029 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301), .A(b_man[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2952));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1030 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2779), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1031 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3445), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1032 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3301), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3102));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1033 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1034 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3716), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1035 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1036 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3581), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1037 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1038 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2246), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1039 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3375), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3240), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3508));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1040 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2248), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3370), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2452));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1041 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2189), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2754), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3425));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1042 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1043 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2417), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1044 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2746), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1045 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1046 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2885), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1047 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2382), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2527));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1048 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2379), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2805), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2678), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3159));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1049 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3227), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3639), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3027));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1050 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3507), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2962), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2333));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1051 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1052 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1053 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1054 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3168), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1055 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1056 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3034), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1057 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028), .A(b_man[5]), .B(b_man[6]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1058 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369), .A(b_man[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3028));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1059 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1060 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3641), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1061 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3369), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3303));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1062 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2813), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2668), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3085));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1063 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2661), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3709), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2609));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1064 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1065 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1066 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2306), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1067 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1068 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2176), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1069 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2453), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2871), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2531), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3228));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1070 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3439), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3710));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1071 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2872), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2512), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2878));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1072 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1073 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1074 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1075 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2956), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1076 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1077 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3096), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1078 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2593), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2741));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1079 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3285), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2725), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3148));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1080 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1081 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090), .A(b_man[3]), .B(b_man[4]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1082 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430), .A(b_man[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3090));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1083 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2988), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1084 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2239), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1085 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3430), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3504));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1086 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1087 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3234), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1088 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3484), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2877), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2934));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1089 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1090 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1091 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2520), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2941), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2377), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3291));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1092 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1093 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2373), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1094 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2624), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1095 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3161), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1096 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1097 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3298), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1098 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2807), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2948));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1099 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2168), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3635), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2788));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1101 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1102 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1103 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154), .A(b_man[1]), .B(b_man[2]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1104 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495), .A(b_man[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3154));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1105 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2268), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2448), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1107 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3495), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3705));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2588), .A1(N13252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2237), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3357));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1110 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3529), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361));
OA22X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3364), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2655), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3361), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2721));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1115 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1116 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1117 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2233), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3342));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1118 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1119 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3695), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3353));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3683), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2426));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1122 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3141), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2220));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3294), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2946));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2574), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3625));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1126 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1127 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2362), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3424));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1128 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1129 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2310), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3577));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2162), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3567));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1131 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1132 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2814));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1133 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2764), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2401));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1135 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3167), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3647));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1136 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1137 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2389), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3253));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3591), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2836));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1140 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2460), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3717));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1141 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3195), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3132));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1142 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3476), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3418));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1143 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446));
AOI31X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1144 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706), .A2(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3231));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1145 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2153), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2444));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1146 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2806), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3100));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1147 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2388), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3649));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1149 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3442), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2828));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3188), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2560));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1152 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2916), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2644));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1154 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3338), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2993));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1155 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3362), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3019));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1156 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739));
AOI2BB2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1157 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3012), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2739), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1158 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3093), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3517));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2257), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2700));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1160 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3314), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2968));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3471), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3646), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3308));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1162 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3064), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2224));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2579), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3374));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1164 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3112), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3656), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2757));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1165 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3714), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2902));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1166 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3257), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3139));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2904), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2546));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2563), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3446), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2384), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3107));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6892 (.Y(N13270), .A(N11981));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6893 (.Y(N13273), .A(N11983), .B(N11829));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6894 (.Y(N13271), .A(N13270), .B(N13273));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6895 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557), .A(N13271));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1170 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3481), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3368));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1171 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3707), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2894));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1172 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2692), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3256), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2331));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1173 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3250), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2777));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3129), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3215));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1175 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2483), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3055), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3740));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3249), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2185), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2893));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1177 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3558), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2375));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1178 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2742), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2468));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1179 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2274), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3537));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2825), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2915));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3266), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2286));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1182 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3680), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3341));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1183 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3050), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2685));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1184 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2651), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2715), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3275), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2350));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1185 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441), .A0(N11973), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557), .B0(N11971));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1186 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2641), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3630));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1187 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2670), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2368));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1188 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3480), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2423), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3138));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1189 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3035), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3660));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1190 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3600));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1191 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3284), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2219), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2930));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1192 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2835), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3389), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2476));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1193 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2334), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2277));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1194 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2634), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3485));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1195 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3082), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3623), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2724));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1196 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2223), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3426));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1197 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2300), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2164));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1198 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2869), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3422), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2509));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1199 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2621), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3191), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2267));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1200 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2501), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3073), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2150));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1201 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3099), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3360));
AOI31X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1202 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440), .A0(N11962), .A1(N11812), .A2(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441), .B0(N11960));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1203 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2663), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3171));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1204 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3312));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1205 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2659), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3225), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2297));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1206 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3652));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1207 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3254), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2900));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2449), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3025), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3708));
OA21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1209 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2342), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2415), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2986), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3672));
OAI31X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1210 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707), .A0(N11951), .A1(N11664), .A2(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440), .B0(N11949));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1211 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2811), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2481), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3594));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1212 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542), .A0(N11319), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707), .B0(N11941));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1213 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3011));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1214 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2977));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1215 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2992), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2838));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6896 (.Y(N13280), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3542), .B(N11930));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6897 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47]), .A(N13280));
INVXL buf1_A_I6907 (.Y(N13319), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47]));
INVXL buf1_A_I6908 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360), .A(N13319));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6876 (.Y(N13253), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6885 (.Y(N13262), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6884 (.Y(N13261), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6883 (.Y(N13260), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6882 (.Y(N13259), .A(N13253));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6881 (.Y(N13258), .A(N13253));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6880 (.Y(N13257), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6879 (.Y(N13256), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6878 (.Y(N13255), .A(N13253));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6877 (.Y(N13254), .A(N13253));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1218 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2707), .B(N11319));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1219 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47]), .A(N13254), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1220 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1221 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336), .A0(N11343), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383), .B0(N11552));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1222 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2336), .B(N11307));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1223 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914), .A0(N11664), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3440), .B0(N11662));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1224 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914), .B(N11325));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1225 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44]), .S0(N13256));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1226 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2383), .B(N11343));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1227 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[43]), .S0(N13254));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1228 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1229 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746), .A0(N11325), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2914), .B0(N11539));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1230 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3746), .B(N11301));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1231 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[46]), .S0(N13255));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1232 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[44]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[45]), .S0(N13255));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1233 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1234 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5506));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1235 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1236 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176), .A0(N11684), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306), .B0(N11717));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1238 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3176), .B(N11536));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325), .A0(N11712), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3163), .B0(N11710));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325), .B(N11549));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36]), .S0(N13257));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1242 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3306), .B(N11684));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[35]), .S0(N13257));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1244 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972), .A0(N11549), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3325), .B0(N11573));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1246 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2972), .B(N11337));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1247 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637), .A0(N11812), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2441), .B0(N11810));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1248 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1249 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643), .B(N11355));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1250 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38]), .S0(N13256));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1251 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2669), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2995));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1252 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2824), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2324));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1253 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157), .A(N12649));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1254 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497), .A(N12652));
OA21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6898 (.Y(N13287), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3157), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3497));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6899 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235), .A(N13287));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3185), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3589));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1257 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522), .A0(N11906), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235), .B0(N11904));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1258 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3036), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2629));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1259 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376), .A0(N11793), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522), .B0(N11791));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1260 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3376), .B(N11658));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1261 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[34]), .S0(N13258));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1262 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3522), .B(N11672));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1263 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[33]), .S0(N13257));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2171), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3197));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1266 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2235));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1267 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2524), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2842));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1268 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879), .A0(N11804), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958), .B0(N11802));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2879), .B(N11678));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1270 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[32]), .S0(N13258));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2958), .B(N11702));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[31]), .S0(N13257));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1273 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5526), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1275 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[37]), .S0(N13254));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1276 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1278 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584), .A0(N11727), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595), .B0(N11742));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2584), .B(N11583));
OA21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6900 (.Y(N13294), .A0(N11758), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3557), .B0(N11756));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6901 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044), .A(N13294));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044), .B(N11589));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28]), .S0(N13257));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1283 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2595), .B(N11727));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1284 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[27]), .S0(N13256));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1285 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367), .A0(N11589), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3044), .B0(N11592));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2367), .B(N11361));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1288 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[30]), .S0(N13256));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1289 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3694), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2193));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1290 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530), .A(N12655));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1291 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886), .A(N12658));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1292 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2530), .A1(N11829), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2886));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1293 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2435), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3454));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1294 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798), .A0(N11823), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242), .B0(N11821));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1295 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2798), .B(N11733));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[26]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3242), .B(N11739));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[25]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1300 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285), .A0(N11831), .A1(N11829), .B0(N11840));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1301 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2285), .B(N11752));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1302 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[24]), .S0(N13258));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1303 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1304 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5547), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1305 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[29]), .S0(N13255));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1306 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1307 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5496), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1308 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121), .A0(N11694), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3637), .B0(N11692));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1309 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550), .A0(N11349), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121), .B0(N11559));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1310 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2550), .B(N11313));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1311 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[42]), .S0(N13255));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1312 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3121), .B(N11349));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1313 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[41]), .S0(N13255));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761), .A0(N11355), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3643), .B0(N11566));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2761), .B(N11331));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1317 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[40]), .S0(N13256));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1318 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[38]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[39]), .S0(N13254));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1319 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1320 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1321 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5473), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1322 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[47]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8442));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1323 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22]), .A(N11829), .B(N11831));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[23]), .S0(N13254));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1326 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1327 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23), .A(a_sign), .B(b_sign));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1328 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N445), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1329 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1330 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1331 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1332 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3678), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3701));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1333 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2782), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3134));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1334 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2738));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1335 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2]), .A(N11465), .B(N11467), .S0(N13259));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1336 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3280), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3621));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1337 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3411), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2672));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1338 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2358), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2719));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1339 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2802), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3722));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1340 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6]), .A(N11453), .B(N11488), .S0(N13259));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3478), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2215));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2830), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2174));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2569), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2928));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2413), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3237));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1345 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4]), .A(N11507), .B(N11451), .S0(N13260));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3080), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3420));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3582), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3179));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2156), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2507));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1349 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2767), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2613));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1350 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8]), .A(N11495), .B(N11472), .S0(N13260));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1351 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[4]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[8]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2866), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3221));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1353 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3349), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3663));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1354 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3118));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10]), .A(N11458), .B(N11460), .S0(N13258));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1358 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2446), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2808));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3169), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3063));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1360 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2491));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1362 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14]), .A(N11479), .B(N11481), .S0(N13259));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2294), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2307));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2209), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3561));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2656), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3022));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1366 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2158), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2553));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1367 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3365), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3706));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1368 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2486), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3603));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1369 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12]), .A(N11500), .B(N11502), .S0(N13260));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1370 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3502), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2247));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1371 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3072), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3162));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1372 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2240), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2594));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1373 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3563), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3546));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1374 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1375 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3005));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1376 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16]), .A(N11521), .B(N11523), .S0(N13260));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1377 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[10]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[14]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[12]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[16]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1378 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5]), .A(N11451), .B(N11453), .S0(N13258));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1379 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9]), .A(N11472), .B(N11458), .S0(N13259));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1380 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7]), .A(N11488), .B(N11495), .S0(N13259));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11]), .A(N11460), .B(N11500), .S0(N13260));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1382 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[9]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[7]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[11]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3]), .A(N11467), .B(N11507), .S0(N13261));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1384 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1385 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2252));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2495), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3405), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3755));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21]), .A(N11835), .B(N11837));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1388 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[22]), .S0(N13262));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1389 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[22]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1390 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2459), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3513));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1391 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2600), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2606));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1392 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20]), .A(N11624), .B(N12644), .S0(N13261));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1393 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3304), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2954));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1394 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3642), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2380));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3669), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2431));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1396 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2155));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1397 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3417));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1398 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3137), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3617), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2784));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1399 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2747), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3103));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1400 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2772), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N3489));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1401 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18]), .A(N11643), .B(N11645), .S0(N13262));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[20]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[18]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[0]), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2293));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0]), .A(N13261), .B(N11610));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1]), .A(N11610), .B(N11465), .S0(N13261));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1406 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21]), .A(N12644), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[21]), .S0(N13261));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1407 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13]), .A(N11502), .B(N11479), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17]), .A(N11523), .B(N11643), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5360));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1409 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15]), .A(N11481), .B(N11521), .S0(N13262));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19]), .A(N11645), .B(N11624), .S0(N13262));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6902 (.Y(N13303), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[13]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[17]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[15]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6903 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679), .A(N13303));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1412 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[1]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[21]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5679));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1413 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5664), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5674), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5692));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1414 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5672), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5662), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5688), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5666));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[24]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N443), .B(N10969), .C(N10971), .D(N10973));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447), .A(N10921), .B(N10923), .C(N10925), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N444));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450), .A0(N10923), .A1(N10925), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__34));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[23]), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N447), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N450));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6904 (.Y(N13309), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__24[47]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6905 (.Y(N13311), .A(N13309));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6906 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38), .A(N13311));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1421 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0]), .A(N10812), .B(N10814), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1422 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1423 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5765));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1425 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5758));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1426 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1427 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]), .A(N10858), .B(N10860), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1428 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5777));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1429 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5831));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1431 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5789));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1432 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1433 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]), .A(N10867), .B(N10869), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1434 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1435 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5771));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1436 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5815), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1437 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]), .A(N10821), .B(N10823), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1438 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1439 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5786));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1440 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[5]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5835));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1441 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1442 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761), .A(a_exp[7]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1443 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5761), .B(b_exp[7]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5766));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5833), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7]), .A(N10876), .B(N10878), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1446 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5816), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[3]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]), .A(N10885), .B(N10887), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1449 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8]), .A(a_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1450 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1451 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8]), .A(N10798), .B(N10800), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5834), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[6]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]), .A(N10830), .B(N10832), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1454 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[1]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1455 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]), .A(N10839), .B(N10841), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1456 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5825));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1457 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9]), .A(a_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5781));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1458 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__31[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5824), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1459 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]), .A(N10790), .B(N10792), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__38));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1460 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]));
NOR3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1461 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5949));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1462 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__20), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__13));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1463 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__21), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__14));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1464 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964), .A(N10751), .B(N10753), .C(N9758), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1465 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5946), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5942), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5964));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1466 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[5]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1467 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[2]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1468 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[3]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1469 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5909), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5897));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1470 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5904));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1471 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5906), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8450));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1472 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N461));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1473 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N8456), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[9]));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1474 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__49), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5957), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__51));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123), .A(N12662));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082), .A(N10567), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6886 (.Y(N13263), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6082));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6887 (.Y(N13264), .A(N13263));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1477 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178), .A(N13264), .B(N10230));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1478 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5502), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1480 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .A(N10645), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123), .B(N10645));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081), .A0(N10422), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10428));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1483 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6144), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192), .A(N10593), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6888 (.Y(N13265), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6192));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6889 (.Y(N13266), .A(N13265));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1485 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106), .A(N10619), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6123));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6890 (.Y(N13267), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6106));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I6891 (.Y(N13268), .A(N13267));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1486 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986), .A(rm[0]), .B(rm[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1487 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7), .A(rm[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5986));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1488 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__7), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__6));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1489 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5634), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__5));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1490 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1491 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[7]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1492 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__30[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N442));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1493 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6044), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1494 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173), .A0(N10114), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1495 (.Y(x[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6081), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6173));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1496 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095), .A(N13264), .B(N10225));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1498 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[44]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191), .A0(N10413), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10419));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199), .A0(N10105), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1501 (.Y(x[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6095), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6191), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6199));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1502 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205), .A(N13264), .B(N10220));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1503 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1504 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5477), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[43]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1505 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107), .A0(N10404), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10410));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1506 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221), .A0(N10096), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1507 (.Y(x[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6205), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6107), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6221));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1508 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120), .A(N13264), .B(N10215));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1509 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1510 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5505), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[42]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1511 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214), .A0(N10395), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10401));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1512 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247), .A0(N10087), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1513 (.Y(x[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6120), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6214), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6247));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228), .A(N13264), .B(N10210));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1515 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5557), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1516 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5540), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[41]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1517 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132), .A0(N10386), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10392));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1518 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078), .A0(N10078), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1519 (.Y(x[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6132), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6078));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1520 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146), .A(N13264), .B(N10205));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1522 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5480), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[40]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239), .A0(N10377), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10383));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1524 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103), .A0(N10069), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1525 (.Y(x[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6146), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6239), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6103));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061), .A(N13264), .B(N10200));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1527 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[39]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1528 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157), .A0(N10368), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10374));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1529 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129), .A0(N10060), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1530 (.Y(x[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6061), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6157), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6129));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168), .A(N13264), .B(N10195));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1533 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5554), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1534 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5530), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[38]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1535 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071), .A0(N10359), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10365));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1536 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154), .A0(N10051), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1537 (.Y(x[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6168), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6071), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6154));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085), .A(N13264), .B(N10190));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1539 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5489), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1540 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5495), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[37]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1541 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181), .A0(N10350), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10356));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1542 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177), .A0(N10042), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1543 (.Y(x[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6085), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6181), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6177));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1544 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193), .A(N13264), .B(N10185));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1545 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1546 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5487), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[36]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097), .A0(N10341), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10347));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1548 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203), .A0(N10033), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1549 (.Y(x[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6193), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6097), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6203));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1550 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110), .A(N13264), .B(N10180));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1551 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5501));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1552 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[35]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1553 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207), .A0(N10332), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10338));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1554 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226), .A0(N10024), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1555 (.Y(x[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6110), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6207), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6226));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1556 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216), .A(N13264), .B(N10175));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1557 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1558 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[34]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1559 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122), .A0(N10323), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10329));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060), .A0(N10015), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1561 (.Y(x[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6216), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6122), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6060));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1562 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135), .A(N13264), .B(N10170));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1563 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5539), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[33]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1565 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230), .A0(N10314), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10320));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083), .A0(N10006), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1567 (.Y(x[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6135), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6230), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6083));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1568 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242), .A(N13264), .B(N10165));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1569 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1570 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5497), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[32]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1571 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148), .A0(N10305), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10311));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108), .A0(N9997), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1573 (.Y(x[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6242), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6148), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6108));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162), .A(N13264), .B(N10160));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1575 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[31]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1576 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063), .A0(N10296), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10302));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1577 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134), .A0(N9988), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1578 (.Y(x[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6162), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6063), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6134));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1579 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073), .A(N13264), .B(N10155));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1581 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5542), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[30]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1582 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170), .A0(N10287), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10293));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1583 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160), .A0(N9979), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1584 (.Y(x[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6073), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6170), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6160));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1585 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185), .A(N13264), .B(N10150));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1586 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1587 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5482), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[29]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1588 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087), .A0(N10278), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10284));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183), .A0(N9970), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1590 (.Y(x[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6185), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6087), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6183));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100), .A(N13264), .B(N10145));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1592 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1593 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[28]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1594 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196), .A0(N10269), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10275));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1595 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209), .A0(N9961), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1596 (.Y(x[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6100), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6196), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6209));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1597 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210), .A(N13264), .B(N10140));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1598 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5523), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[27]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1599 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112), .A0(N10260), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10266));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1600 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232), .A0(N9952), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1601 (.Y(x[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6210), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6112), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6232));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1602 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126), .A(N13264), .B(N10135));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1603 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1604 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5474), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[26]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1605 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218), .A0(N10251), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10257));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1606 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064), .A0(N9943), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1607 (.Y(x[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6126), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6218), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6064));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1608 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234), .A(N13264), .B(N10130));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1609 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[25]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1610 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138), .A0(N10242), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10248));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1611 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089), .A0(N9934), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1612 (.Y(x[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6234), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6138), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6089));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1613 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150), .A(N13264), .B(N10125));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1614 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244), .A0(N10233), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6158), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6117), .B1(N10239));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1615 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114), .A0(N9925), .A1(N13266), .B0(N13268), .B1(N13250));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1616 (.Y(x[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6150), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6244), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6114));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1617 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5507), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[45]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5528), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5520));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1618 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N5472), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1619 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6053), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__25[46]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__44));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1620 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__47));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1621 (.Y(x[22]), .A(N9680), .B(N9678), .S0(N13248));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1622 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__32));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1623 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__27), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1624 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6008), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1625 (.Y(x[30]), .A(N9624), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1626 (.Y(x[29]), .A(N9631), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1627 (.Y(x[28]), .A(N9638), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1628 (.Y(x[27]), .A(N9645), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1629 (.Y(x[26]), .A(N9652), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1630 (.Y(x[25]), .A(N9659), .B(N9633), .S0(N13248));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1631 (.Y(x[24]), .A(N9666), .B(N9633), .S0(N13248));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1632 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6004), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__48[0]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1633 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N6025), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__42), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N469), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N470));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1634 (.Y(x[23]), .A(N9673), .B(N9671), .S0(N13248));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1635 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131), .AN(b_sign), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1636 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2131), .B(a_sign), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__15));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_5_I1637 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__23), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_N2136), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__26));
reg x_reg_L0_31__I1669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I1669_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[31];
	end
assign N4120 = x_reg_L0_31__I1669_QOUT;
reg x_reg_L1_31__I1701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1701_QOUT <= N4120;
	end
assign x[31] = x_reg_L1_31__I1701_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_3_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vLP3Tg3arxo= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



