/****************************************************************************
*
*  Copyright (c) 2015, Cadence Design Systems. All Rights Reserved.
*
*  This file contains confidential information that may not be
*  distributed under any circumstances without the written permision
*  of Cadence Design Systems.
*
****************************************************************************/
/****************************************************************************
*
* Verilog Verification wrapper module for the cache module.
*
* This module contains the followng items:
*	- A foreign module definition for use in instantiatin the type_wrapper module
*      which contains the BEH module instance.
*	- An instance of the type_wrapper foreign module.
*   - alwyas blocks each type_wrapper output.
*
****************************************************************************/

`timescale 1 ps / 1 ps

module cache_vlwrapper(
      clk,
       rstn,
       cache_en,
       systolic_en,
       systolic_depth,
       addr_if_start,
       systolic_sel,
       feature_data,
       feature_share_en,
       feature_data_en,
       feature_data_sel,
       weight_data,
       weight_data_en,
       mac_src_0_s0_0,
      mac_src_0_s0_1,
      mac_src_0_s0_2,
      mac_src_0_s0_3,
      mac_src_0_s0_4,
      mac_src_0_s0_5,
      mac_src_0_s0_6,
      mac_src_0_s0_7,
      mac_src_0_s0_8,
      mac_src_0_s0_9,
      mac_src_0_s0_10,
      mac_src_0_s0_11,
      mac_src_0_s0_12,
      mac_src_0_s0_13,
      mac_src_0_s0_14,
      mac_src_0_s0_15,
      mac_src_0_s0_16,
      mac_src_0_s0_17,
      mac_src_0_s0_18,
      mac_src_0_s0_19,
      mac_src_0_s0_20,
      mac_src_0_s0_21,
      mac_src_0_s0_22,
      mac_src_0_s0_23,
      mac_src_0_s0_24,
      mac_src_0_s0_25,
      mac_src_0_s0_26,
      mac_src_0_s0_27,
      mac_src_0_s0_28,
      mac_src_0_s0_29,
      mac_src_0_s0_30,
      mac_src_0_s0_31,
       mac_src_0_s1_0,
      mac_src_0_s1_1,
      mac_src_0_s1_2,
      mac_src_0_s1_3,
      mac_src_0_s1_4,
      mac_src_0_s1_5,
      mac_src_0_s1_6,
      mac_src_0_s1_7,
      mac_src_0_s1_8,
      mac_src_0_s1_9,
      mac_src_0_s1_10,
      mac_src_0_s1_11,
      mac_src_0_s1_12,
      mac_src_0_s1_13,
      mac_src_0_s1_14,
      mac_src_0_s1_15,
      mac_src_0_s1_16,
      mac_src_0_s1_17,
      mac_src_0_s1_18,
      mac_src_0_s1_19,
      mac_src_0_s1_20,
      mac_src_0_s1_21,
      mac_src_0_s1_22,
      mac_src_0_s1_23,
      mac_src_0_s1_24,
      mac_src_0_s1_25,
      mac_src_0_s1_26,
      mac_src_0_s1_27,
      mac_src_0_s1_28,
      mac_src_0_s1_29,
      mac_src_0_s1_30,
      mac_src_0_s1_31,
       mac_src_0_s2_0,
      mac_src_0_s2_1,
      mac_src_0_s2_2,
      mac_src_0_s2_3,
      mac_src_0_s2_4,
      mac_src_0_s2_5,
      mac_src_0_s2_6,
      mac_src_0_s2_7,
      mac_src_0_s2_8,
      mac_src_0_s2_9,
      mac_src_0_s2_10,
      mac_src_0_s2_11,
      mac_src_0_s2_12,
      mac_src_0_s2_13,
      mac_src_0_s2_14,
      mac_src_0_s2_15,
      mac_src_0_s2_16,
      mac_src_0_s2_17,
      mac_src_0_s2_18,
      mac_src_0_s2_19,
      mac_src_0_s2_20,
      mac_src_0_s2_21,
      mac_src_0_s2_22,
      mac_src_0_s2_23,
      mac_src_0_s2_24,
      mac_src_0_s2_25,
      mac_src_0_s2_26,
      mac_src_0_s2_27,
      mac_src_0_s2_28,
      mac_src_0_s2_29,
      mac_src_0_s2_30,
      mac_src_0_s2_31,
       mac_src_0_s3_0,
      mac_src_0_s3_1,
      mac_src_0_s3_2,
      mac_src_0_s3_3,
      mac_src_0_s3_4,
      mac_src_0_s3_5,
      mac_src_0_s3_6,
      mac_src_0_s3_7,
      mac_src_0_s3_8,
      mac_src_0_s3_9,
      mac_src_0_s3_10,
      mac_src_0_s3_11,
      mac_src_0_s3_12,
      mac_src_0_s3_13,
      mac_src_0_s3_14,
      mac_src_0_s3_15,
      mac_src_0_s3_16,
      mac_src_0_s3_17,
      mac_src_0_s3_18,
      mac_src_0_s3_19,
      mac_src_0_s3_20,
      mac_src_0_s3_21,
      mac_src_0_s3_22,
      mac_src_0_s3_23,
      mac_src_0_s3_24,
      mac_src_0_s3_25,
      mac_src_0_s3_26,
      mac_src_0_s3_27,
      mac_src_0_s3_28,
      mac_src_0_s3_29,
      mac_src_0_s3_30,
      mac_src_0_s3_31,
       mac_src_0_s4_0,
      mac_src_0_s4_1,
      mac_src_0_s4_2,
      mac_src_0_s4_3,
      mac_src_0_s4_4,
      mac_src_0_s4_5,
      mac_src_0_s4_6,
      mac_src_0_s4_7,
      mac_src_0_s4_8,
      mac_src_0_s4_9,
      mac_src_0_s4_10,
      mac_src_0_s4_11,
      mac_src_0_s4_12,
      mac_src_0_s4_13,
      mac_src_0_s4_14,
      mac_src_0_s4_15,
      mac_src_0_s4_16,
      mac_src_0_s4_17,
      mac_src_0_s4_18,
      mac_src_0_s4_19,
      mac_src_0_s4_20,
      mac_src_0_s4_21,
      mac_src_0_s4_22,
      mac_src_0_s4_23,
      mac_src_0_s4_24,
      mac_src_0_s4_25,
      mac_src_0_s4_26,
      mac_src_0_s4_27,
      mac_src_0_s4_28,
      mac_src_0_s4_29,
      mac_src_0_s4_30,
      mac_src_0_s4_31,
       mac_src_0_s5_0,
      mac_src_0_s5_1,
      mac_src_0_s5_2,
      mac_src_0_s5_3,
      mac_src_0_s5_4,
      mac_src_0_s5_5,
      mac_src_0_s5_6,
      mac_src_0_s5_7,
      mac_src_0_s5_8,
      mac_src_0_s5_9,
      mac_src_0_s5_10,
      mac_src_0_s5_11,
      mac_src_0_s5_12,
      mac_src_0_s5_13,
      mac_src_0_s5_14,
      mac_src_0_s5_15,
      mac_src_0_s5_16,
      mac_src_0_s5_17,
      mac_src_0_s5_18,
      mac_src_0_s5_19,
      mac_src_0_s5_20,
      mac_src_0_s5_21,
      mac_src_0_s5_22,
      mac_src_0_s5_23,
      mac_src_0_s5_24,
      mac_src_0_s5_25,
      mac_src_0_s5_26,
      mac_src_0_s5_27,
      mac_src_0_s5_28,
      mac_src_0_s5_29,
      mac_src_0_s5_30,
      mac_src_0_s5_31,
       mac_src_0_s6_0,
      mac_src_0_s6_1,
      mac_src_0_s6_2,
      mac_src_0_s6_3,
      mac_src_0_s6_4,
      mac_src_0_s6_5,
      mac_src_0_s6_6,
      mac_src_0_s6_7,
      mac_src_0_s6_8,
      mac_src_0_s6_9,
      mac_src_0_s6_10,
      mac_src_0_s6_11,
      mac_src_0_s6_12,
      mac_src_0_s6_13,
      mac_src_0_s6_14,
      mac_src_0_s6_15,
      mac_src_0_s6_16,
      mac_src_0_s6_17,
      mac_src_0_s6_18,
      mac_src_0_s6_19,
      mac_src_0_s6_20,
      mac_src_0_s6_21,
      mac_src_0_s6_22,
      mac_src_0_s6_23,
      mac_src_0_s6_24,
      mac_src_0_s6_25,
      mac_src_0_s6_26,
      mac_src_0_s6_27,
      mac_src_0_s6_28,
      mac_src_0_s6_29,
      mac_src_0_s6_30,
      mac_src_0_s6_31,
       mac_src_1_0,
      mac_src_1_1,
      mac_src_1_2,
      mac_src_1_3,
      mac_src_1_4,
      mac_src_1_5,
      mac_src_1_6,
      mac_src_1_7,
      mac_src_1_8,
      mac_src_1_9,
      mac_src_1_10,
      mac_src_1_11,
      mac_src_1_12,
      mac_src_1_13,
      mac_src_1_14,
      mac_src_1_15,
      mac_src_1_16,
      mac_src_1_17,
      mac_src_1_18,
      mac_src_1_19,
      mac_src_1_20,
      mac_src_1_21,
      mac_src_1_22,
      mac_src_1_23,
      mac_src_1_24,
      mac_src_1_25,
      mac_src_1_26,
      mac_src_1_27,
      mac_src_1_28,
      mac_src_1_29,
      mac_src_1_30,
      mac_src_1_31,
       mac_src_valid,
       mac_clear

    );

	input clk;
	input rstn;
	input cache_en;
	input [7:0] systolic_en;
	input [7:0] systolic_depth;
	input addr_if_start;
	input [7:0] systolic_sel;
	input [319:0] feature_data;
	input feature_share_en;
	input feature_data_en;
	input [15:0] feature_data_sel;
	input [255:0] weight_data;
	input weight_data_en;
	output [9:0] mac_src_0_s0_0;
	output [9:0] mac_src_0_s0_1;
	output [9:0] mac_src_0_s0_2;
	output [9:0] mac_src_0_s0_3;
	output [9:0] mac_src_0_s0_4;
	output [9:0] mac_src_0_s0_5;
	output [9:0] mac_src_0_s0_6;
	output [9:0] mac_src_0_s0_7;
	output [9:0] mac_src_0_s0_8;
	output [9:0] mac_src_0_s0_9;
	output [9:0] mac_src_0_s0_10;
	output [9:0] mac_src_0_s0_11;
	output [9:0] mac_src_0_s0_12;
	output [9:0] mac_src_0_s0_13;
	output [9:0] mac_src_0_s0_14;
	output [9:0] mac_src_0_s0_15;
	output [9:0] mac_src_0_s0_16;
	output [9:0] mac_src_0_s0_17;
	output [9:0] mac_src_0_s0_18;
	output [9:0] mac_src_0_s0_19;
	output [9:0] mac_src_0_s0_20;
	output [9:0] mac_src_0_s0_21;
	output [9:0] mac_src_0_s0_22;
	output [9:0] mac_src_0_s0_23;
	output [9:0] mac_src_0_s0_24;
	output [9:0] mac_src_0_s0_25;
	output [9:0] mac_src_0_s0_26;
	output [9:0] mac_src_0_s0_27;
	output [9:0] mac_src_0_s0_28;
	output [9:0] mac_src_0_s0_29;
	output [9:0] mac_src_0_s0_30;
	output [9:0] mac_src_0_s0_31;
	reg[9:0] mac_src_0_s0_0;
	wire [9:0] m_mac_src_0_s0_0;
	reg[9:0] mac_src_0_s0_1;
	wire [9:0] m_mac_src_0_s0_1;
	reg[9:0] mac_src_0_s0_2;
	wire [9:0] m_mac_src_0_s0_2;
	reg[9:0] mac_src_0_s0_3;
	wire [9:0] m_mac_src_0_s0_3;
	reg[9:0] mac_src_0_s0_4;
	wire [9:0] m_mac_src_0_s0_4;
	reg[9:0] mac_src_0_s0_5;
	wire [9:0] m_mac_src_0_s0_5;
	reg[9:0] mac_src_0_s0_6;
	wire [9:0] m_mac_src_0_s0_6;
	reg[9:0] mac_src_0_s0_7;
	wire [9:0] m_mac_src_0_s0_7;
	reg[9:0] mac_src_0_s0_8;
	wire [9:0] m_mac_src_0_s0_8;
	reg[9:0] mac_src_0_s0_9;
	wire [9:0] m_mac_src_0_s0_9;
	reg[9:0] mac_src_0_s0_10;
	wire [9:0] m_mac_src_0_s0_10;
	reg[9:0] mac_src_0_s0_11;
	wire [9:0] m_mac_src_0_s0_11;
	reg[9:0] mac_src_0_s0_12;
	wire [9:0] m_mac_src_0_s0_12;
	reg[9:0] mac_src_0_s0_13;
	wire [9:0] m_mac_src_0_s0_13;
	reg[9:0] mac_src_0_s0_14;
	wire [9:0] m_mac_src_0_s0_14;
	reg[9:0] mac_src_0_s0_15;
	wire [9:0] m_mac_src_0_s0_15;
	reg[9:0] mac_src_0_s0_16;
	wire [9:0] m_mac_src_0_s0_16;
	reg[9:0] mac_src_0_s0_17;
	wire [9:0] m_mac_src_0_s0_17;
	reg[9:0] mac_src_0_s0_18;
	wire [9:0] m_mac_src_0_s0_18;
	reg[9:0] mac_src_0_s0_19;
	wire [9:0] m_mac_src_0_s0_19;
	reg[9:0] mac_src_0_s0_20;
	wire [9:0] m_mac_src_0_s0_20;
	reg[9:0] mac_src_0_s0_21;
	wire [9:0] m_mac_src_0_s0_21;
	reg[9:0] mac_src_0_s0_22;
	wire [9:0] m_mac_src_0_s0_22;
	reg[9:0] mac_src_0_s0_23;
	wire [9:0] m_mac_src_0_s0_23;
	reg[9:0] mac_src_0_s0_24;
	wire [9:0] m_mac_src_0_s0_24;
	reg[9:0] mac_src_0_s0_25;
	wire [9:0] m_mac_src_0_s0_25;
	reg[9:0] mac_src_0_s0_26;
	wire [9:0] m_mac_src_0_s0_26;
	reg[9:0] mac_src_0_s0_27;
	wire [9:0] m_mac_src_0_s0_27;
	reg[9:0] mac_src_0_s0_28;
	wire [9:0] m_mac_src_0_s0_28;
	reg[9:0] mac_src_0_s0_29;
	wire [9:0] m_mac_src_0_s0_29;
	reg[9:0] mac_src_0_s0_30;
	wire [9:0] m_mac_src_0_s0_30;
	reg[9:0] mac_src_0_s0_31;
	wire [9:0] m_mac_src_0_s0_31;
	output [9:0] mac_src_0_s1_0;
	output [9:0] mac_src_0_s1_1;
	output [9:0] mac_src_0_s1_2;
	output [9:0] mac_src_0_s1_3;
	output [9:0] mac_src_0_s1_4;
	output [9:0] mac_src_0_s1_5;
	output [9:0] mac_src_0_s1_6;
	output [9:0] mac_src_0_s1_7;
	output [9:0] mac_src_0_s1_8;
	output [9:0] mac_src_0_s1_9;
	output [9:0] mac_src_0_s1_10;
	output [9:0] mac_src_0_s1_11;
	output [9:0] mac_src_0_s1_12;
	output [9:0] mac_src_0_s1_13;
	output [9:0] mac_src_0_s1_14;
	output [9:0] mac_src_0_s1_15;
	output [9:0] mac_src_0_s1_16;
	output [9:0] mac_src_0_s1_17;
	output [9:0] mac_src_0_s1_18;
	output [9:0] mac_src_0_s1_19;
	output [9:0] mac_src_0_s1_20;
	output [9:0] mac_src_0_s1_21;
	output [9:0] mac_src_0_s1_22;
	output [9:0] mac_src_0_s1_23;
	output [9:0] mac_src_0_s1_24;
	output [9:0] mac_src_0_s1_25;
	output [9:0] mac_src_0_s1_26;
	output [9:0] mac_src_0_s1_27;
	output [9:0] mac_src_0_s1_28;
	output [9:0] mac_src_0_s1_29;
	output [9:0] mac_src_0_s1_30;
	output [9:0] mac_src_0_s1_31;
	reg[9:0] mac_src_0_s1_0;
	wire [9:0] m_mac_src_0_s1_0;
	reg[9:0] mac_src_0_s1_1;
	wire [9:0] m_mac_src_0_s1_1;
	reg[9:0] mac_src_0_s1_2;
	wire [9:0] m_mac_src_0_s1_2;
	reg[9:0] mac_src_0_s1_3;
	wire [9:0] m_mac_src_0_s1_3;
	reg[9:0] mac_src_0_s1_4;
	wire [9:0] m_mac_src_0_s1_4;
	reg[9:0] mac_src_0_s1_5;
	wire [9:0] m_mac_src_0_s1_5;
	reg[9:0] mac_src_0_s1_6;
	wire [9:0] m_mac_src_0_s1_6;
	reg[9:0] mac_src_0_s1_7;
	wire [9:0] m_mac_src_0_s1_7;
	reg[9:0] mac_src_0_s1_8;
	wire [9:0] m_mac_src_0_s1_8;
	reg[9:0] mac_src_0_s1_9;
	wire [9:0] m_mac_src_0_s1_9;
	reg[9:0] mac_src_0_s1_10;
	wire [9:0] m_mac_src_0_s1_10;
	reg[9:0] mac_src_0_s1_11;
	wire [9:0] m_mac_src_0_s1_11;
	reg[9:0] mac_src_0_s1_12;
	wire [9:0] m_mac_src_0_s1_12;
	reg[9:0] mac_src_0_s1_13;
	wire [9:0] m_mac_src_0_s1_13;
	reg[9:0] mac_src_0_s1_14;
	wire [9:0] m_mac_src_0_s1_14;
	reg[9:0] mac_src_0_s1_15;
	wire [9:0] m_mac_src_0_s1_15;
	reg[9:0] mac_src_0_s1_16;
	wire [9:0] m_mac_src_0_s1_16;
	reg[9:0] mac_src_0_s1_17;
	wire [9:0] m_mac_src_0_s1_17;
	reg[9:0] mac_src_0_s1_18;
	wire [9:0] m_mac_src_0_s1_18;
	reg[9:0] mac_src_0_s1_19;
	wire [9:0] m_mac_src_0_s1_19;
	reg[9:0] mac_src_0_s1_20;
	wire [9:0] m_mac_src_0_s1_20;
	reg[9:0] mac_src_0_s1_21;
	wire [9:0] m_mac_src_0_s1_21;
	reg[9:0] mac_src_0_s1_22;
	wire [9:0] m_mac_src_0_s1_22;
	reg[9:0] mac_src_0_s1_23;
	wire [9:0] m_mac_src_0_s1_23;
	reg[9:0] mac_src_0_s1_24;
	wire [9:0] m_mac_src_0_s1_24;
	reg[9:0] mac_src_0_s1_25;
	wire [9:0] m_mac_src_0_s1_25;
	reg[9:0] mac_src_0_s1_26;
	wire [9:0] m_mac_src_0_s1_26;
	reg[9:0] mac_src_0_s1_27;
	wire [9:0] m_mac_src_0_s1_27;
	reg[9:0] mac_src_0_s1_28;
	wire [9:0] m_mac_src_0_s1_28;
	reg[9:0] mac_src_0_s1_29;
	wire [9:0] m_mac_src_0_s1_29;
	reg[9:0] mac_src_0_s1_30;
	wire [9:0] m_mac_src_0_s1_30;
	reg[9:0] mac_src_0_s1_31;
	wire [9:0] m_mac_src_0_s1_31;
	output [9:0] mac_src_0_s2_0;
	output [9:0] mac_src_0_s2_1;
	output [9:0] mac_src_0_s2_2;
	output [9:0] mac_src_0_s2_3;
	output [9:0] mac_src_0_s2_4;
	output [9:0] mac_src_0_s2_5;
	output [9:0] mac_src_0_s2_6;
	output [9:0] mac_src_0_s2_7;
	output [9:0] mac_src_0_s2_8;
	output [9:0] mac_src_0_s2_9;
	output [9:0] mac_src_0_s2_10;
	output [9:0] mac_src_0_s2_11;
	output [9:0] mac_src_0_s2_12;
	output [9:0] mac_src_0_s2_13;
	output [9:0] mac_src_0_s2_14;
	output [9:0] mac_src_0_s2_15;
	output [9:0] mac_src_0_s2_16;
	output [9:0] mac_src_0_s2_17;
	output [9:0] mac_src_0_s2_18;
	output [9:0] mac_src_0_s2_19;
	output [9:0] mac_src_0_s2_20;
	output [9:0] mac_src_0_s2_21;
	output [9:0] mac_src_0_s2_22;
	output [9:0] mac_src_0_s2_23;
	output [9:0] mac_src_0_s2_24;
	output [9:0] mac_src_0_s2_25;
	output [9:0] mac_src_0_s2_26;
	output [9:0] mac_src_0_s2_27;
	output [9:0] mac_src_0_s2_28;
	output [9:0] mac_src_0_s2_29;
	output [9:0] mac_src_0_s2_30;
	output [9:0] mac_src_0_s2_31;
	reg[9:0] mac_src_0_s2_0;
	wire [9:0] m_mac_src_0_s2_0;
	reg[9:0] mac_src_0_s2_1;
	wire [9:0] m_mac_src_0_s2_1;
	reg[9:0] mac_src_0_s2_2;
	wire [9:0] m_mac_src_0_s2_2;
	reg[9:0] mac_src_0_s2_3;
	wire [9:0] m_mac_src_0_s2_3;
	reg[9:0] mac_src_0_s2_4;
	wire [9:0] m_mac_src_0_s2_4;
	reg[9:0] mac_src_0_s2_5;
	wire [9:0] m_mac_src_0_s2_5;
	reg[9:0] mac_src_0_s2_6;
	wire [9:0] m_mac_src_0_s2_6;
	reg[9:0] mac_src_0_s2_7;
	wire [9:0] m_mac_src_0_s2_7;
	reg[9:0] mac_src_0_s2_8;
	wire [9:0] m_mac_src_0_s2_8;
	reg[9:0] mac_src_0_s2_9;
	wire [9:0] m_mac_src_0_s2_9;
	reg[9:0] mac_src_0_s2_10;
	wire [9:0] m_mac_src_0_s2_10;
	reg[9:0] mac_src_0_s2_11;
	wire [9:0] m_mac_src_0_s2_11;
	reg[9:0] mac_src_0_s2_12;
	wire [9:0] m_mac_src_0_s2_12;
	reg[9:0] mac_src_0_s2_13;
	wire [9:0] m_mac_src_0_s2_13;
	reg[9:0] mac_src_0_s2_14;
	wire [9:0] m_mac_src_0_s2_14;
	reg[9:0] mac_src_0_s2_15;
	wire [9:0] m_mac_src_0_s2_15;
	reg[9:0] mac_src_0_s2_16;
	wire [9:0] m_mac_src_0_s2_16;
	reg[9:0] mac_src_0_s2_17;
	wire [9:0] m_mac_src_0_s2_17;
	reg[9:0] mac_src_0_s2_18;
	wire [9:0] m_mac_src_0_s2_18;
	reg[9:0] mac_src_0_s2_19;
	wire [9:0] m_mac_src_0_s2_19;
	reg[9:0] mac_src_0_s2_20;
	wire [9:0] m_mac_src_0_s2_20;
	reg[9:0] mac_src_0_s2_21;
	wire [9:0] m_mac_src_0_s2_21;
	reg[9:0] mac_src_0_s2_22;
	wire [9:0] m_mac_src_0_s2_22;
	reg[9:0] mac_src_0_s2_23;
	wire [9:0] m_mac_src_0_s2_23;
	reg[9:0] mac_src_0_s2_24;
	wire [9:0] m_mac_src_0_s2_24;
	reg[9:0] mac_src_0_s2_25;
	wire [9:0] m_mac_src_0_s2_25;
	reg[9:0] mac_src_0_s2_26;
	wire [9:0] m_mac_src_0_s2_26;
	reg[9:0] mac_src_0_s2_27;
	wire [9:0] m_mac_src_0_s2_27;
	reg[9:0] mac_src_0_s2_28;
	wire [9:0] m_mac_src_0_s2_28;
	reg[9:0] mac_src_0_s2_29;
	wire [9:0] m_mac_src_0_s2_29;
	reg[9:0] mac_src_0_s2_30;
	wire [9:0] m_mac_src_0_s2_30;
	reg[9:0] mac_src_0_s2_31;
	wire [9:0] m_mac_src_0_s2_31;
	output [9:0] mac_src_0_s3_0;
	output [9:0] mac_src_0_s3_1;
	output [9:0] mac_src_0_s3_2;
	output [9:0] mac_src_0_s3_3;
	output [9:0] mac_src_0_s3_4;
	output [9:0] mac_src_0_s3_5;
	output [9:0] mac_src_0_s3_6;
	output [9:0] mac_src_0_s3_7;
	output [9:0] mac_src_0_s3_8;
	output [9:0] mac_src_0_s3_9;
	output [9:0] mac_src_0_s3_10;
	output [9:0] mac_src_0_s3_11;
	output [9:0] mac_src_0_s3_12;
	output [9:0] mac_src_0_s3_13;
	output [9:0] mac_src_0_s3_14;
	output [9:0] mac_src_0_s3_15;
	output [9:0] mac_src_0_s3_16;
	output [9:0] mac_src_0_s3_17;
	output [9:0] mac_src_0_s3_18;
	output [9:0] mac_src_0_s3_19;
	output [9:0] mac_src_0_s3_20;
	output [9:0] mac_src_0_s3_21;
	output [9:0] mac_src_0_s3_22;
	output [9:0] mac_src_0_s3_23;
	output [9:0] mac_src_0_s3_24;
	output [9:0] mac_src_0_s3_25;
	output [9:0] mac_src_0_s3_26;
	output [9:0] mac_src_0_s3_27;
	output [9:0] mac_src_0_s3_28;
	output [9:0] mac_src_0_s3_29;
	output [9:0] mac_src_0_s3_30;
	output [9:0] mac_src_0_s3_31;
	reg[9:0] mac_src_0_s3_0;
	wire [9:0] m_mac_src_0_s3_0;
	reg[9:0] mac_src_0_s3_1;
	wire [9:0] m_mac_src_0_s3_1;
	reg[9:0] mac_src_0_s3_2;
	wire [9:0] m_mac_src_0_s3_2;
	reg[9:0] mac_src_0_s3_3;
	wire [9:0] m_mac_src_0_s3_3;
	reg[9:0] mac_src_0_s3_4;
	wire [9:0] m_mac_src_0_s3_4;
	reg[9:0] mac_src_0_s3_5;
	wire [9:0] m_mac_src_0_s3_5;
	reg[9:0] mac_src_0_s3_6;
	wire [9:0] m_mac_src_0_s3_6;
	reg[9:0] mac_src_0_s3_7;
	wire [9:0] m_mac_src_0_s3_7;
	reg[9:0] mac_src_0_s3_8;
	wire [9:0] m_mac_src_0_s3_8;
	reg[9:0] mac_src_0_s3_9;
	wire [9:0] m_mac_src_0_s3_9;
	reg[9:0] mac_src_0_s3_10;
	wire [9:0] m_mac_src_0_s3_10;
	reg[9:0] mac_src_0_s3_11;
	wire [9:0] m_mac_src_0_s3_11;
	reg[9:0] mac_src_0_s3_12;
	wire [9:0] m_mac_src_0_s3_12;
	reg[9:0] mac_src_0_s3_13;
	wire [9:0] m_mac_src_0_s3_13;
	reg[9:0] mac_src_0_s3_14;
	wire [9:0] m_mac_src_0_s3_14;
	reg[9:0] mac_src_0_s3_15;
	wire [9:0] m_mac_src_0_s3_15;
	reg[9:0] mac_src_0_s3_16;
	wire [9:0] m_mac_src_0_s3_16;
	reg[9:0] mac_src_0_s3_17;
	wire [9:0] m_mac_src_0_s3_17;
	reg[9:0] mac_src_0_s3_18;
	wire [9:0] m_mac_src_0_s3_18;
	reg[9:0] mac_src_0_s3_19;
	wire [9:0] m_mac_src_0_s3_19;
	reg[9:0] mac_src_0_s3_20;
	wire [9:0] m_mac_src_0_s3_20;
	reg[9:0] mac_src_0_s3_21;
	wire [9:0] m_mac_src_0_s3_21;
	reg[9:0] mac_src_0_s3_22;
	wire [9:0] m_mac_src_0_s3_22;
	reg[9:0] mac_src_0_s3_23;
	wire [9:0] m_mac_src_0_s3_23;
	reg[9:0] mac_src_0_s3_24;
	wire [9:0] m_mac_src_0_s3_24;
	reg[9:0] mac_src_0_s3_25;
	wire [9:0] m_mac_src_0_s3_25;
	reg[9:0] mac_src_0_s3_26;
	wire [9:0] m_mac_src_0_s3_26;
	reg[9:0] mac_src_0_s3_27;
	wire [9:0] m_mac_src_0_s3_27;
	reg[9:0] mac_src_0_s3_28;
	wire [9:0] m_mac_src_0_s3_28;
	reg[9:0] mac_src_0_s3_29;
	wire [9:0] m_mac_src_0_s3_29;
	reg[9:0] mac_src_0_s3_30;
	wire [9:0] m_mac_src_0_s3_30;
	reg[9:0] mac_src_0_s3_31;
	wire [9:0] m_mac_src_0_s3_31;
	output [9:0] mac_src_0_s4_0;
	output [9:0] mac_src_0_s4_1;
	output [9:0] mac_src_0_s4_2;
	output [9:0] mac_src_0_s4_3;
	output [9:0] mac_src_0_s4_4;
	output [9:0] mac_src_0_s4_5;
	output [9:0] mac_src_0_s4_6;
	output [9:0] mac_src_0_s4_7;
	output [9:0] mac_src_0_s4_8;
	output [9:0] mac_src_0_s4_9;
	output [9:0] mac_src_0_s4_10;
	output [9:0] mac_src_0_s4_11;
	output [9:0] mac_src_0_s4_12;
	output [9:0] mac_src_0_s4_13;
	output [9:0] mac_src_0_s4_14;
	output [9:0] mac_src_0_s4_15;
	output [9:0] mac_src_0_s4_16;
	output [9:0] mac_src_0_s4_17;
	output [9:0] mac_src_0_s4_18;
	output [9:0] mac_src_0_s4_19;
	output [9:0] mac_src_0_s4_20;
	output [9:0] mac_src_0_s4_21;
	output [9:0] mac_src_0_s4_22;
	output [9:0] mac_src_0_s4_23;
	output [9:0] mac_src_0_s4_24;
	output [9:0] mac_src_0_s4_25;
	output [9:0] mac_src_0_s4_26;
	output [9:0] mac_src_0_s4_27;
	output [9:0] mac_src_0_s4_28;
	output [9:0] mac_src_0_s4_29;
	output [9:0] mac_src_0_s4_30;
	output [9:0] mac_src_0_s4_31;
	reg[9:0] mac_src_0_s4_0;
	wire [9:0] m_mac_src_0_s4_0;
	reg[9:0] mac_src_0_s4_1;
	wire [9:0] m_mac_src_0_s4_1;
	reg[9:0] mac_src_0_s4_2;
	wire [9:0] m_mac_src_0_s4_2;
	reg[9:0] mac_src_0_s4_3;
	wire [9:0] m_mac_src_0_s4_3;
	reg[9:0] mac_src_0_s4_4;
	wire [9:0] m_mac_src_0_s4_4;
	reg[9:0] mac_src_0_s4_5;
	wire [9:0] m_mac_src_0_s4_5;
	reg[9:0] mac_src_0_s4_6;
	wire [9:0] m_mac_src_0_s4_6;
	reg[9:0] mac_src_0_s4_7;
	wire [9:0] m_mac_src_0_s4_7;
	reg[9:0] mac_src_0_s4_8;
	wire [9:0] m_mac_src_0_s4_8;
	reg[9:0] mac_src_0_s4_9;
	wire [9:0] m_mac_src_0_s4_9;
	reg[9:0] mac_src_0_s4_10;
	wire [9:0] m_mac_src_0_s4_10;
	reg[9:0] mac_src_0_s4_11;
	wire [9:0] m_mac_src_0_s4_11;
	reg[9:0] mac_src_0_s4_12;
	wire [9:0] m_mac_src_0_s4_12;
	reg[9:0] mac_src_0_s4_13;
	wire [9:0] m_mac_src_0_s4_13;
	reg[9:0] mac_src_0_s4_14;
	wire [9:0] m_mac_src_0_s4_14;
	reg[9:0] mac_src_0_s4_15;
	wire [9:0] m_mac_src_0_s4_15;
	reg[9:0] mac_src_0_s4_16;
	wire [9:0] m_mac_src_0_s4_16;
	reg[9:0] mac_src_0_s4_17;
	wire [9:0] m_mac_src_0_s4_17;
	reg[9:0] mac_src_0_s4_18;
	wire [9:0] m_mac_src_0_s4_18;
	reg[9:0] mac_src_0_s4_19;
	wire [9:0] m_mac_src_0_s4_19;
	reg[9:0] mac_src_0_s4_20;
	wire [9:0] m_mac_src_0_s4_20;
	reg[9:0] mac_src_0_s4_21;
	wire [9:0] m_mac_src_0_s4_21;
	reg[9:0] mac_src_0_s4_22;
	wire [9:0] m_mac_src_0_s4_22;
	reg[9:0] mac_src_0_s4_23;
	wire [9:0] m_mac_src_0_s4_23;
	reg[9:0] mac_src_0_s4_24;
	wire [9:0] m_mac_src_0_s4_24;
	reg[9:0] mac_src_0_s4_25;
	wire [9:0] m_mac_src_0_s4_25;
	reg[9:0] mac_src_0_s4_26;
	wire [9:0] m_mac_src_0_s4_26;
	reg[9:0] mac_src_0_s4_27;
	wire [9:0] m_mac_src_0_s4_27;
	reg[9:0] mac_src_0_s4_28;
	wire [9:0] m_mac_src_0_s4_28;
	reg[9:0] mac_src_0_s4_29;
	wire [9:0] m_mac_src_0_s4_29;
	reg[9:0] mac_src_0_s4_30;
	wire [9:0] m_mac_src_0_s4_30;
	reg[9:0] mac_src_0_s4_31;
	wire [9:0] m_mac_src_0_s4_31;
	output [9:0] mac_src_0_s5_0;
	output [9:0] mac_src_0_s5_1;
	output [9:0] mac_src_0_s5_2;
	output [9:0] mac_src_0_s5_3;
	output [9:0] mac_src_0_s5_4;
	output [9:0] mac_src_0_s5_5;
	output [9:0] mac_src_0_s5_6;
	output [9:0] mac_src_0_s5_7;
	output [9:0] mac_src_0_s5_8;
	output [9:0] mac_src_0_s5_9;
	output [9:0] mac_src_0_s5_10;
	output [9:0] mac_src_0_s5_11;
	output [9:0] mac_src_0_s5_12;
	output [9:0] mac_src_0_s5_13;
	output [9:0] mac_src_0_s5_14;
	output [9:0] mac_src_0_s5_15;
	output [9:0] mac_src_0_s5_16;
	output [9:0] mac_src_0_s5_17;
	output [9:0] mac_src_0_s5_18;
	output [9:0] mac_src_0_s5_19;
	output [9:0] mac_src_0_s5_20;
	output [9:0] mac_src_0_s5_21;
	output [9:0] mac_src_0_s5_22;
	output [9:0] mac_src_0_s5_23;
	output [9:0] mac_src_0_s5_24;
	output [9:0] mac_src_0_s5_25;
	output [9:0] mac_src_0_s5_26;
	output [9:0] mac_src_0_s5_27;
	output [9:0] mac_src_0_s5_28;
	output [9:0] mac_src_0_s5_29;
	output [9:0] mac_src_0_s5_30;
	output [9:0] mac_src_0_s5_31;
	reg[9:0] mac_src_0_s5_0;
	wire [9:0] m_mac_src_0_s5_0;
	reg[9:0] mac_src_0_s5_1;
	wire [9:0] m_mac_src_0_s5_1;
	reg[9:0] mac_src_0_s5_2;
	wire [9:0] m_mac_src_0_s5_2;
	reg[9:0] mac_src_0_s5_3;
	wire [9:0] m_mac_src_0_s5_3;
	reg[9:0] mac_src_0_s5_4;
	wire [9:0] m_mac_src_0_s5_4;
	reg[9:0] mac_src_0_s5_5;
	wire [9:0] m_mac_src_0_s5_5;
	reg[9:0] mac_src_0_s5_6;
	wire [9:0] m_mac_src_0_s5_6;
	reg[9:0] mac_src_0_s5_7;
	wire [9:0] m_mac_src_0_s5_7;
	reg[9:0] mac_src_0_s5_8;
	wire [9:0] m_mac_src_0_s5_8;
	reg[9:0] mac_src_0_s5_9;
	wire [9:0] m_mac_src_0_s5_9;
	reg[9:0] mac_src_0_s5_10;
	wire [9:0] m_mac_src_0_s5_10;
	reg[9:0] mac_src_0_s5_11;
	wire [9:0] m_mac_src_0_s5_11;
	reg[9:0] mac_src_0_s5_12;
	wire [9:0] m_mac_src_0_s5_12;
	reg[9:0] mac_src_0_s5_13;
	wire [9:0] m_mac_src_0_s5_13;
	reg[9:0] mac_src_0_s5_14;
	wire [9:0] m_mac_src_0_s5_14;
	reg[9:0] mac_src_0_s5_15;
	wire [9:0] m_mac_src_0_s5_15;
	reg[9:0] mac_src_0_s5_16;
	wire [9:0] m_mac_src_0_s5_16;
	reg[9:0] mac_src_0_s5_17;
	wire [9:0] m_mac_src_0_s5_17;
	reg[9:0] mac_src_0_s5_18;
	wire [9:0] m_mac_src_0_s5_18;
	reg[9:0] mac_src_0_s5_19;
	wire [9:0] m_mac_src_0_s5_19;
	reg[9:0] mac_src_0_s5_20;
	wire [9:0] m_mac_src_0_s5_20;
	reg[9:0] mac_src_0_s5_21;
	wire [9:0] m_mac_src_0_s5_21;
	reg[9:0] mac_src_0_s5_22;
	wire [9:0] m_mac_src_0_s5_22;
	reg[9:0] mac_src_0_s5_23;
	wire [9:0] m_mac_src_0_s5_23;
	reg[9:0] mac_src_0_s5_24;
	wire [9:0] m_mac_src_0_s5_24;
	reg[9:0] mac_src_0_s5_25;
	wire [9:0] m_mac_src_0_s5_25;
	reg[9:0] mac_src_0_s5_26;
	wire [9:0] m_mac_src_0_s5_26;
	reg[9:0] mac_src_0_s5_27;
	wire [9:0] m_mac_src_0_s5_27;
	reg[9:0] mac_src_0_s5_28;
	wire [9:0] m_mac_src_0_s5_28;
	reg[9:0] mac_src_0_s5_29;
	wire [9:0] m_mac_src_0_s5_29;
	reg[9:0] mac_src_0_s5_30;
	wire [9:0] m_mac_src_0_s5_30;
	reg[9:0] mac_src_0_s5_31;
	wire [9:0] m_mac_src_0_s5_31;
	output [9:0] mac_src_0_s6_0;
	output [9:0] mac_src_0_s6_1;
	output [9:0] mac_src_0_s6_2;
	output [9:0] mac_src_0_s6_3;
	output [9:0] mac_src_0_s6_4;
	output [9:0] mac_src_0_s6_5;
	output [9:0] mac_src_0_s6_6;
	output [9:0] mac_src_0_s6_7;
	output [9:0] mac_src_0_s6_8;
	output [9:0] mac_src_0_s6_9;
	output [9:0] mac_src_0_s6_10;
	output [9:0] mac_src_0_s6_11;
	output [9:0] mac_src_0_s6_12;
	output [9:0] mac_src_0_s6_13;
	output [9:0] mac_src_0_s6_14;
	output [9:0] mac_src_0_s6_15;
	output [9:0] mac_src_0_s6_16;
	output [9:0] mac_src_0_s6_17;
	output [9:0] mac_src_0_s6_18;
	output [9:0] mac_src_0_s6_19;
	output [9:0] mac_src_0_s6_20;
	output [9:0] mac_src_0_s6_21;
	output [9:0] mac_src_0_s6_22;
	output [9:0] mac_src_0_s6_23;
	output [9:0] mac_src_0_s6_24;
	output [9:0] mac_src_0_s6_25;
	output [9:0] mac_src_0_s6_26;
	output [9:0] mac_src_0_s6_27;
	output [9:0] mac_src_0_s6_28;
	output [9:0] mac_src_0_s6_29;
	output [9:0] mac_src_0_s6_30;
	output [9:0] mac_src_0_s6_31;
	reg[9:0] mac_src_0_s6_0;
	wire [9:0] m_mac_src_0_s6_0;
	reg[9:0] mac_src_0_s6_1;
	wire [9:0] m_mac_src_0_s6_1;
	reg[9:0] mac_src_0_s6_2;
	wire [9:0] m_mac_src_0_s6_2;
	reg[9:0] mac_src_0_s6_3;
	wire [9:0] m_mac_src_0_s6_3;
	reg[9:0] mac_src_0_s6_4;
	wire [9:0] m_mac_src_0_s6_4;
	reg[9:0] mac_src_0_s6_5;
	wire [9:0] m_mac_src_0_s6_5;
	reg[9:0] mac_src_0_s6_6;
	wire [9:0] m_mac_src_0_s6_6;
	reg[9:0] mac_src_0_s6_7;
	wire [9:0] m_mac_src_0_s6_7;
	reg[9:0] mac_src_0_s6_8;
	wire [9:0] m_mac_src_0_s6_8;
	reg[9:0] mac_src_0_s6_9;
	wire [9:0] m_mac_src_0_s6_9;
	reg[9:0] mac_src_0_s6_10;
	wire [9:0] m_mac_src_0_s6_10;
	reg[9:0] mac_src_0_s6_11;
	wire [9:0] m_mac_src_0_s6_11;
	reg[9:0] mac_src_0_s6_12;
	wire [9:0] m_mac_src_0_s6_12;
	reg[9:0] mac_src_0_s6_13;
	wire [9:0] m_mac_src_0_s6_13;
	reg[9:0] mac_src_0_s6_14;
	wire [9:0] m_mac_src_0_s6_14;
	reg[9:0] mac_src_0_s6_15;
	wire [9:0] m_mac_src_0_s6_15;
	reg[9:0] mac_src_0_s6_16;
	wire [9:0] m_mac_src_0_s6_16;
	reg[9:0] mac_src_0_s6_17;
	wire [9:0] m_mac_src_0_s6_17;
	reg[9:0] mac_src_0_s6_18;
	wire [9:0] m_mac_src_0_s6_18;
	reg[9:0] mac_src_0_s6_19;
	wire [9:0] m_mac_src_0_s6_19;
	reg[9:0] mac_src_0_s6_20;
	wire [9:0] m_mac_src_0_s6_20;
	reg[9:0] mac_src_0_s6_21;
	wire [9:0] m_mac_src_0_s6_21;
	reg[9:0] mac_src_0_s6_22;
	wire [9:0] m_mac_src_0_s6_22;
	reg[9:0] mac_src_0_s6_23;
	wire [9:0] m_mac_src_0_s6_23;
	reg[9:0] mac_src_0_s6_24;
	wire [9:0] m_mac_src_0_s6_24;
	reg[9:0] mac_src_0_s6_25;
	wire [9:0] m_mac_src_0_s6_25;
	reg[9:0] mac_src_0_s6_26;
	wire [9:0] m_mac_src_0_s6_26;
	reg[9:0] mac_src_0_s6_27;
	wire [9:0] m_mac_src_0_s6_27;
	reg[9:0] mac_src_0_s6_28;
	wire [9:0] m_mac_src_0_s6_28;
	reg[9:0] mac_src_0_s6_29;
	wire [9:0] m_mac_src_0_s6_29;
	reg[9:0] mac_src_0_s6_30;
	wire [9:0] m_mac_src_0_s6_30;
	reg[9:0] mac_src_0_s6_31;
	wire [9:0] m_mac_src_0_s6_31;
	output [7:0] mac_src_1_0;
	output [7:0] mac_src_1_1;
	output [7:0] mac_src_1_2;
	output [7:0] mac_src_1_3;
	output [7:0] mac_src_1_4;
	output [7:0] mac_src_1_5;
	output [7:0] mac_src_1_6;
	output [7:0] mac_src_1_7;
	output [7:0] mac_src_1_8;
	output [7:0] mac_src_1_9;
	output [7:0] mac_src_1_10;
	output [7:0] mac_src_1_11;
	output [7:0] mac_src_1_12;
	output [7:0] mac_src_1_13;
	output [7:0] mac_src_1_14;
	output [7:0] mac_src_1_15;
	output [7:0] mac_src_1_16;
	output [7:0] mac_src_1_17;
	output [7:0] mac_src_1_18;
	output [7:0] mac_src_1_19;
	output [7:0] mac_src_1_20;
	output [7:0] mac_src_1_21;
	output [7:0] mac_src_1_22;
	output [7:0] mac_src_1_23;
	output [7:0] mac_src_1_24;
	output [7:0] mac_src_1_25;
	output [7:0] mac_src_1_26;
	output [7:0] mac_src_1_27;
	output [7:0] mac_src_1_28;
	output [7:0] mac_src_1_29;
	output [7:0] mac_src_1_30;
	output [7:0] mac_src_1_31;
	reg[7:0] mac_src_1_0;
	wire [7:0] m_mac_src_1_0;
	reg[7:0] mac_src_1_1;
	wire [7:0] m_mac_src_1_1;
	reg[7:0] mac_src_1_2;
	wire [7:0] m_mac_src_1_2;
	reg[7:0] mac_src_1_3;
	wire [7:0] m_mac_src_1_3;
	reg[7:0] mac_src_1_4;
	wire [7:0] m_mac_src_1_4;
	reg[7:0] mac_src_1_5;
	wire [7:0] m_mac_src_1_5;
	reg[7:0] mac_src_1_6;
	wire [7:0] m_mac_src_1_6;
	reg[7:0] mac_src_1_7;
	wire [7:0] m_mac_src_1_7;
	reg[7:0] mac_src_1_8;
	wire [7:0] m_mac_src_1_8;
	reg[7:0] mac_src_1_9;
	wire [7:0] m_mac_src_1_9;
	reg[7:0] mac_src_1_10;
	wire [7:0] m_mac_src_1_10;
	reg[7:0] mac_src_1_11;
	wire [7:0] m_mac_src_1_11;
	reg[7:0] mac_src_1_12;
	wire [7:0] m_mac_src_1_12;
	reg[7:0] mac_src_1_13;
	wire [7:0] m_mac_src_1_13;
	reg[7:0] mac_src_1_14;
	wire [7:0] m_mac_src_1_14;
	reg[7:0] mac_src_1_15;
	wire [7:0] m_mac_src_1_15;
	reg[7:0] mac_src_1_16;
	wire [7:0] m_mac_src_1_16;
	reg[7:0] mac_src_1_17;
	wire [7:0] m_mac_src_1_17;
	reg[7:0] mac_src_1_18;
	wire [7:0] m_mac_src_1_18;
	reg[7:0] mac_src_1_19;
	wire [7:0] m_mac_src_1_19;
	reg[7:0] mac_src_1_20;
	wire [7:0] m_mac_src_1_20;
	reg[7:0] mac_src_1_21;
	wire [7:0] m_mac_src_1_21;
	reg[7:0] mac_src_1_22;
	wire [7:0] m_mac_src_1_22;
	reg[7:0] mac_src_1_23;
	wire [7:0] m_mac_src_1_23;
	reg[7:0] mac_src_1_24;
	wire [7:0] m_mac_src_1_24;
	reg[7:0] mac_src_1_25;
	wire [7:0] m_mac_src_1_25;
	reg[7:0] mac_src_1_26;
	wire [7:0] m_mac_src_1_26;
	reg[7:0] mac_src_1_27;
	wire [7:0] m_mac_src_1_27;
	reg[7:0] mac_src_1_28;
	wire [7:0] m_mac_src_1_28;
	reg[7:0] mac_src_1_29;
	wire [7:0] m_mac_src_1_29;
	reg[7:0] mac_src_1_30;
	wire [7:0] m_mac_src_1_30;
	reg[7:0] mac_src_1_31;
	wire [7:0] m_mac_src_1_31;
	output mac_src_valid;
	reg mac_src_valid;
	wire m_mac_src_valid;
	output mac_clear;
	reg mac_clear;
	wire m_mac_clear;


    // Instantiate the Verilog module that instantiates the SystemC module
    cache_type_wrapper cache_sc(
        .clk(clk),
         .rstn(rstn),
         .cache_en(cache_en),
         .systolic_en(systolic_en),
         .systolic_depth(systolic_depth),
         .addr_if_start(addr_if_start),
         .systolic_sel(systolic_sel),
         .feature_data(feature_data),
         .feature_share_en(feature_share_en),
         .feature_data_en(feature_data_en),
         .feature_data_sel(feature_data_sel),
         .weight_data(weight_data),
         .weight_data_en(weight_data_en),
         .mac_src_0_s0_0(m_mac_src_0_s0_0),
        .mac_src_0_s0_1(m_mac_src_0_s0_1),
        .mac_src_0_s0_2(m_mac_src_0_s0_2),
        .mac_src_0_s0_3(m_mac_src_0_s0_3),
        .mac_src_0_s0_4(m_mac_src_0_s0_4),
        .mac_src_0_s0_5(m_mac_src_0_s0_5),
        .mac_src_0_s0_6(m_mac_src_0_s0_6),
        .mac_src_0_s0_7(m_mac_src_0_s0_7),
        .mac_src_0_s0_8(m_mac_src_0_s0_8),
        .mac_src_0_s0_9(m_mac_src_0_s0_9),
        .mac_src_0_s0_10(m_mac_src_0_s0_10),
        .mac_src_0_s0_11(m_mac_src_0_s0_11),
        .mac_src_0_s0_12(m_mac_src_0_s0_12),
        .mac_src_0_s0_13(m_mac_src_0_s0_13),
        .mac_src_0_s0_14(m_mac_src_0_s0_14),
        .mac_src_0_s0_15(m_mac_src_0_s0_15),
        .mac_src_0_s0_16(m_mac_src_0_s0_16),
        .mac_src_0_s0_17(m_mac_src_0_s0_17),
        .mac_src_0_s0_18(m_mac_src_0_s0_18),
        .mac_src_0_s0_19(m_mac_src_0_s0_19),
        .mac_src_0_s0_20(m_mac_src_0_s0_20),
        .mac_src_0_s0_21(m_mac_src_0_s0_21),
        .mac_src_0_s0_22(m_mac_src_0_s0_22),
        .mac_src_0_s0_23(m_mac_src_0_s0_23),
        .mac_src_0_s0_24(m_mac_src_0_s0_24),
        .mac_src_0_s0_25(m_mac_src_0_s0_25),
        .mac_src_0_s0_26(m_mac_src_0_s0_26),
        .mac_src_0_s0_27(m_mac_src_0_s0_27),
        .mac_src_0_s0_28(m_mac_src_0_s0_28),
        .mac_src_0_s0_29(m_mac_src_0_s0_29),
        .mac_src_0_s0_30(m_mac_src_0_s0_30),
        .mac_src_0_s0_31(m_mac_src_0_s0_31),
         .mac_src_0_s1_0(m_mac_src_0_s1_0),
        .mac_src_0_s1_1(m_mac_src_0_s1_1),
        .mac_src_0_s1_2(m_mac_src_0_s1_2),
        .mac_src_0_s1_3(m_mac_src_0_s1_3),
        .mac_src_0_s1_4(m_mac_src_0_s1_4),
        .mac_src_0_s1_5(m_mac_src_0_s1_5),
        .mac_src_0_s1_6(m_mac_src_0_s1_6),
        .mac_src_0_s1_7(m_mac_src_0_s1_7),
        .mac_src_0_s1_8(m_mac_src_0_s1_8),
        .mac_src_0_s1_9(m_mac_src_0_s1_9),
        .mac_src_0_s1_10(m_mac_src_0_s1_10),
        .mac_src_0_s1_11(m_mac_src_0_s1_11),
        .mac_src_0_s1_12(m_mac_src_0_s1_12),
        .mac_src_0_s1_13(m_mac_src_0_s1_13),
        .mac_src_0_s1_14(m_mac_src_0_s1_14),
        .mac_src_0_s1_15(m_mac_src_0_s1_15),
        .mac_src_0_s1_16(m_mac_src_0_s1_16),
        .mac_src_0_s1_17(m_mac_src_0_s1_17),
        .mac_src_0_s1_18(m_mac_src_0_s1_18),
        .mac_src_0_s1_19(m_mac_src_0_s1_19),
        .mac_src_0_s1_20(m_mac_src_0_s1_20),
        .mac_src_0_s1_21(m_mac_src_0_s1_21),
        .mac_src_0_s1_22(m_mac_src_0_s1_22),
        .mac_src_0_s1_23(m_mac_src_0_s1_23),
        .mac_src_0_s1_24(m_mac_src_0_s1_24),
        .mac_src_0_s1_25(m_mac_src_0_s1_25),
        .mac_src_0_s1_26(m_mac_src_0_s1_26),
        .mac_src_0_s1_27(m_mac_src_0_s1_27),
        .mac_src_0_s1_28(m_mac_src_0_s1_28),
        .mac_src_0_s1_29(m_mac_src_0_s1_29),
        .mac_src_0_s1_30(m_mac_src_0_s1_30),
        .mac_src_0_s1_31(m_mac_src_0_s1_31),
         .mac_src_0_s2_0(m_mac_src_0_s2_0),
        .mac_src_0_s2_1(m_mac_src_0_s2_1),
        .mac_src_0_s2_2(m_mac_src_0_s2_2),
        .mac_src_0_s2_3(m_mac_src_0_s2_3),
        .mac_src_0_s2_4(m_mac_src_0_s2_4),
        .mac_src_0_s2_5(m_mac_src_0_s2_5),
        .mac_src_0_s2_6(m_mac_src_0_s2_6),
        .mac_src_0_s2_7(m_mac_src_0_s2_7),
        .mac_src_0_s2_8(m_mac_src_0_s2_8),
        .mac_src_0_s2_9(m_mac_src_0_s2_9),
        .mac_src_0_s2_10(m_mac_src_0_s2_10),
        .mac_src_0_s2_11(m_mac_src_0_s2_11),
        .mac_src_0_s2_12(m_mac_src_0_s2_12),
        .mac_src_0_s2_13(m_mac_src_0_s2_13),
        .mac_src_0_s2_14(m_mac_src_0_s2_14),
        .mac_src_0_s2_15(m_mac_src_0_s2_15),
        .mac_src_0_s2_16(m_mac_src_0_s2_16),
        .mac_src_0_s2_17(m_mac_src_0_s2_17),
        .mac_src_0_s2_18(m_mac_src_0_s2_18),
        .mac_src_0_s2_19(m_mac_src_0_s2_19),
        .mac_src_0_s2_20(m_mac_src_0_s2_20),
        .mac_src_0_s2_21(m_mac_src_0_s2_21),
        .mac_src_0_s2_22(m_mac_src_0_s2_22),
        .mac_src_0_s2_23(m_mac_src_0_s2_23),
        .mac_src_0_s2_24(m_mac_src_0_s2_24),
        .mac_src_0_s2_25(m_mac_src_0_s2_25),
        .mac_src_0_s2_26(m_mac_src_0_s2_26),
        .mac_src_0_s2_27(m_mac_src_0_s2_27),
        .mac_src_0_s2_28(m_mac_src_0_s2_28),
        .mac_src_0_s2_29(m_mac_src_0_s2_29),
        .mac_src_0_s2_30(m_mac_src_0_s2_30),
        .mac_src_0_s2_31(m_mac_src_0_s2_31),
         .mac_src_0_s3_0(m_mac_src_0_s3_0),
        .mac_src_0_s3_1(m_mac_src_0_s3_1),
        .mac_src_0_s3_2(m_mac_src_0_s3_2),
        .mac_src_0_s3_3(m_mac_src_0_s3_3),
        .mac_src_0_s3_4(m_mac_src_0_s3_4),
        .mac_src_0_s3_5(m_mac_src_0_s3_5),
        .mac_src_0_s3_6(m_mac_src_0_s3_6),
        .mac_src_0_s3_7(m_mac_src_0_s3_7),
        .mac_src_0_s3_8(m_mac_src_0_s3_8),
        .mac_src_0_s3_9(m_mac_src_0_s3_9),
        .mac_src_0_s3_10(m_mac_src_0_s3_10),
        .mac_src_0_s3_11(m_mac_src_0_s3_11),
        .mac_src_0_s3_12(m_mac_src_0_s3_12),
        .mac_src_0_s3_13(m_mac_src_0_s3_13),
        .mac_src_0_s3_14(m_mac_src_0_s3_14),
        .mac_src_0_s3_15(m_mac_src_0_s3_15),
        .mac_src_0_s3_16(m_mac_src_0_s3_16),
        .mac_src_0_s3_17(m_mac_src_0_s3_17),
        .mac_src_0_s3_18(m_mac_src_0_s3_18),
        .mac_src_0_s3_19(m_mac_src_0_s3_19),
        .mac_src_0_s3_20(m_mac_src_0_s3_20),
        .mac_src_0_s3_21(m_mac_src_0_s3_21),
        .mac_src_0_s3_22(m_mac_src_0_s3_22),
        .mac_src_0_s3_23(m_mac_src_0_s3_23),
        .mac_src_0_s3_24(m_mac_src_0_s3_24),
        .mac_src_0_s3_25(m_mac_src_0_s3_25),
        .mac_src_0_s3_26(m_mac_src_0_s3_26),
        .mac_src_0_s3_27(m_mac_src_0_s3_27),
        .mac_src_0_s3_28(m_mac_src_0_s3_28),
        .mac_src_0_s3_29(m_mac_src_0_s3_29),
        .mac_src_0_s3_30(m_mac_src_0_s3_30),
        .mac_src_0_s3_31(m_mac_src_0_s3_31),
         .mac_src_0_s4_0(m_mac_src_0_s4_0),
        .mac_src_0_s4_1(m_mac_src_0_s4_1),
        .mac_src_0_s4_2(m_mac_src_0_s4_2),
        .mac_src_0_s4_3(m_mac_src_0_s4_3),
        .mac_src_0_s4_4(m_mac_src_0_s4_4),
        .mac_src_0_s4_5(m_mac_src_0_s4_5),
        .mac_src_0_s4_6(m_mac_src_0_s4_6),
        .mac_src_0_s4_7(m_mac_src_0_s4_7),
        .mac_src_0_s4_8(m_mac_src_0_s4_8),
        .mac_src_0_s4_9(m_mac_src_0_s4_9),
        .mac_src_0_s4_10(m_mac_src_0_s4_10),
        .mac_src_0_s4_11(m_mac_src_0_s4_11),
        .mac_src_0_s4_12(m_mac_src_0_s4_12),
        .mac_src_0_s4_13(m_mac_src_0_s4_13),
        .mac_src_0_s4_14(m_mac_src_0_s4_14),
        .mac_src_0_s4_15(m_mac_src_0_s4_15),
        .mac_src_0_s4_16(m_mac_src_0_s4_16),
        .mac_src_0_s4_17(m_mac_src_0_s4_17),
        .mac_src_0_s4_18(m_mac_src_0_s4_18),
        .mac_src_0_s4_19(m_mac_src_0_s4_19),
        .mac_src_0_s4_20(m_mac_src_0_s4_20),
        .mac_src_0_s4_21(m_mac_src_0_s4_21),
        .mac_src_0_s4_22(m_mac_src_0_s4_22),
        .mac_src_0_s4_23(m_mac_src_0_s4_23),
        .mac_src_0_s4_24(m_mac_src_0_s4_24),
        .mac_src_0_s4_25(m_mac_src_0_s4_25),
        .mac_src_0_s4_26(m_mac_src_0_s4_26),
        .mac_src_0_s4_27(m_mac_src_0_s4_27),
        .mac_src_0_s4_28(m_mac_src_0_s4_28),
        .mac_src_0_s4_29(m_mac_src_0_s4_29),
        .mac_src_0_s4_30(m_mac_src_0_s4_30),
        .mac_src_0_s4_31(m_mac_src_0_s4_31),
         .mac_src_0_s5_0(m_mac_src_0_s5_0),
        .mac_src_0_s5_1(m_mac_src_0_s5_1),
        .mac_src_0_s5_2(m_mac_src_0_s5_2),
        .mac_src_0_s5_3(m_mac_src_0_s5_3),
        .mac_src_0_s5_4(m_mac_src_0_s5_4),
        .mac_src_0_s5_5(m_mac_src_0_s5_5),
        .mac_src_0_s5_6(m_mac_src_0_s5_6),
        .mac_src_0_s5_7(m_mac_src_0_s5_7),
        .mac_src_0_s5_8(m_mac_src_0_s5_8),
        .mac_src_0_s5_9(m_mac_src_0_s5_9),
        .mac_src_0_s5_10(m_mac_src_0_s5_10),
        .mac_src_0_s5_11(m_mac_src_0_s5_11),
        .mac_src_0_s5_12(m_mac_src_0_s5_12),
        .mac_src_0_s5_13(m_mac_src_0_s5_13),
        .mac_src_0_s5_14(m_mac_src_0_s5_14),
        .mac_src_0_s5_15(m_mac_src_0_s5_15),
        .mac_src_0_s5_16(m_mac_src_0_s5_16),
        .mac_src_0_s5_17(m_mac_src_0_s5_17),
        .mac_src_0_s5_18(m_mac_src_0_s5_18),
        .mac_src_0_s5_19(m_mac_src_0_s5_19),
        .mac_src_0_s5_20(m_mac_src_0_s5_20),
        .mac_src_0_s5_21(m_mac_src_0_s5_21),
        .mac_src_0_s5_22(m_mac_src_0_s5_22),
        .mac_src_0_s5_23(m_mac_src_0_s5_23),
        .mac_src_0_s5_24(m_mac_src_0_s5_24),
        .mac_src_0_s5_25(m_mac_src_0_s5_25),
        .mac_src_0_s5_26(m_mac_src_0_s5_26),
        .mac_src_0_s5_27(m_mac_src_0_s5_27),
        .mac_src_0_s5_28(m_mac_src_0_s5_28),
        .mac_src_0_s5_29(m_mac_src_0_s5_29),
        .mac_src_0_s5_30(m_mac_src_0_s5_30),
        .mac_src_0_s5_31(m_mac_src_0_s5_31),
         .mac_src_0_s6_0(m_mac_src_0_s6_0),
        .mac_src_0_s6_1(m_mac_src_0_s6_1),
        .mac_src_0_s6_2(m_mac_src_0_s6_2),
        .mac_src_0_s6_3(m_mac_src_0_s6_3),
        .mac_src_0_s6_4(m_mac_src_0_s6_4),
        .mac_src_0_s6_5(m_mac_src_0_s6_5),
        .mac_src_0_s6_6(m_mac_src_0_s6_6),
        .mac_src_0_s6_7(m_mac_src_0_s6_7),
        .mac_src_0_s6_8(m_mac_src_0_s6_8),
        .mac_src_0_s6_9(m_mac_src_0_s6_9),
        .mac_src_0_s6_10(m_mac_src_0_s6_10),
        .mac_src_0_s6_11(m_mac_src_0_s6_11),
        .mac_src_0_s6_12(m_mac_src_0_s6_12),
        .mac_src_0_s6_13(m_mac_src_0_s6_13),
        .mac_src_0_s6_14(m_mac_src_0_s6_14),
        .mac_src_0_s6_15(m_mac_src_0_s6_15),
        .mac_src_0_s6_16(m_mac_src_0_s6_16),
        .mac_src_0_s6_17(m_mac_src_0_s6_17),
        .mac_src_0_s6_18(m_mac_src_0_s6_18),
        .mac_src_0_s6_19(m_mac_src_0_s6_19),
        .mac_src_0_s6_20(m_mac_src_0_s6_20),
        .mac_src_0_s6_21(m_mac_src_0_s6_21),
        .mac_src_0_s6_22(m_mac_src_0_s6_22),
        .mac_src_0_s6_23(m_mac_src_0_s6_23),
        .mac_src_0_s6_24(m_mac_src_0_s6_24),
        .mac_src_0_s6_25(m_mac_src_0_s6_25),
        .mac_src_0_s6_26(m_mac_src_0_s6_26),
        .mac_src_0_s6_27(m_mac_src_0_s6_27),
        .mac_src_0_s6_28(m_mac_src_0_s6_28),
        .mac_src_0_s6_29(m_mac_src_0_s6_29),
        .mac_src_0_s6_30(m_mac_src_0_s6_30),
        .mac_src_0_s6_31(m_mac_src_0_s6_31),
         .mac_src_1_0(m_mac_src_1_0),
        .mac_src_1_1(m_mac_src_1_1),
        .mac_src_1_2(m_mac_src_1_2),
        .mac_src_1_3(m_mac_src_1_3),
        .mac_src_1_4(m_mac_src_1_4),
        .mac_src_1_5(m_mac_src_1_5),
        .mac_src_1_6(m_mac_src_1_6),
        .mac_src_1_7(m_mac_src_1_7),
        .mac_src_1_8(m_mac_src_1_8),
        .mac_src_1_9(m_mac_src_1_9),
        .mac_src_1_10(m_mac_src_1_10),
        .mac_src_1_11(m_mac_src_1_11),
        .mac_src_1_12(m_mac_src_1_12),
        .mac_src_1_13(m_mac_src_1_13),
        .mac_src_1_14(m_mac_src_1_14),
        .mac_src_1_15(m_mac_src_1_15),
        .mac_src_1_16(m_mac_src_1_16),
        .mac_src_1_17(m_mac_src_1_17),
        .mac_src_1_18(m_mac_src_1_18),
        .mac_src_1_19(m_mac_src_1_19),
        .mac_src_1_20(m_mac_src_1_20),
        .mac_src_1_21(m_mac_src_1_21),
        .mac_src_1_22(m_mac_src_1_22),
        .mac_src_1_23(m_mac_src_1_23),
        .mac_src_1_24(m_mac_src_1_24),
        .mac_src_1_25(m_mac_src_1_25),
        .mac_src_1_26(m_mac_src_1_26),
        .mac_src_1_27(m_mac_src_1_27),
        .mac_src_1_28(m_mac_src_1_28),
        .mac_src_1_29(m_mac_src_1_29),
        .mac_src_1_30(m_mac_src_1_30),
        .mac_src_1_31(m_mac_src_1_31),
         .mac_src_valid(m_mac_src_valid),
         .mac_clear(m_mac_clear)

    );

    // Always blocks for non-blocking assignments of type_wrapper outputs to
    // Verilog Verificatoin wrapper outputs.

    always @(m_mac_src_0_s0_0)
     begin
      mac_src_0_s0_0 <= m_mac_src_0_s0_0;
     end
    always @(m_mac_src_0_s0_1)
     begin
      mac_src_0_s0_1 <= m_mac_src_0_s0_1;
     end
    always @(m_mac_src_0_s0_2)
     begin
      mac_src_0_s0_2 <= m_mac_src_0_s0_2;
     end
    always @(m_mac_src_0_s0_3)
     begin
      mac_src_0_s0_3 <= m_mac_src_0_s0_3;
     end
    always @(m_mac_src_0_s0_4)
     begin
      mac_src_0_s0_4 <= m_mac_src_0_s0_4;
     end
    always @(m_mac_src_0_s0_5)
     begin
      mac_src_0_s0_5 <= m_mac_src_0_s0_5;
     end
    always @(m_mac_src_0_s0_6)
     begin
      mac_src_0_s0_6 <= m_mac_src_0_s0_6;
     end
    always @(m_mac_src_0_s0_7)
     begin
      mac_src_0_s0_7 <= m_mac_src_0_s0_7;
     end
    always @(m_mac_src_0_s0_8)
     begin
      mac_src_0_s0_8 <= m_mac_src_0_s0_8;
     end
    always @(m_mac_src_0_s0_9)
     begin
      mac_src_0_s0_9 <= m_mac_src_0_s0_9;
     end
    always @(m_mac_src_0_s0_10)
     begin
      mac_src_0_s0_10 <= m_mac_src_0_s0_10;
     end
    always @(m_mac_src_0_s0_11)
     begin
      mac_src_0_s0_11 <= m_mac_src_0_s0_11;
     end
    always @(m_mac_src_0_s0_12)
     begin
      mac_src_0_s0_12 <= m_mac_src_0_s0_12;
     end
    always @(m_mac_src_0_s0_13)
     begin
      mac_src_0_s0_13 <= m_mac_src_0_s0_13;
     end
    always @(m_mac_src_0_s0_14)
     begin
      mac_src_0_s0_14 <= m_mac_src_0_s0_14;
     end
    always @(m_mac_src_0_s0_15)
     begin
      mac_src_0_s0_15 <= m_mac_src_0_s0_15;
     end
    always @(m_mac_src_0_s0_16)
     begin
      mac_src_0_s0_16 <= m_mac_src_0_s0_16;
     end
    always @(m_mac_src_0_s0_17)
     begin
      mac_src_0_s0_17 <= m_mac_src_0_s0_17;
     end
    always @(m_mac_src_0_s0_18)
     begin
      mac_src_0_s0_18 <= m_mac_src_0_s0_18;
     end
    always @(m_mac_src_0_s0_19)
     begin
      mac_src_0_s0_19 <= m_mac_src_0_s0_19;
     end
    always @(m_mac_src_0_s0_20)
     begin
      mac_src_0_s0_20 <= m_mac_src_0_s0_20;
     end
    always @(m_mac_src_0_s0_21)
     begin
      mac_src_0_s0_21 <= m_mac_src_0_s0_21;
     end
    always @(m_mac_src_0_s0_22)
     begin
      mac_src_0_s0_22 <= m_mac_src_0_s0_22;
     end
    always @(m_mac_src_0_s0_23)
     begin
      mac_src_0_s0_23 <= m_mac_src_0_s0_23;
     end
    always @(m_mac_src_0_s0_24)
     begin
      mac_src_0_s0_24 <= m_mac_src_0_s0_24;
     end
    always @(m_mac_src_0_s0_25)
     begin
      mac_src_0_s0_25 <= m_mac_src_0_s0_25;
     end
    always @(m_mac_src_0_s0_26)
     begin
      mac_src_0_s0_26 <= m_mac_src_0_s0_26;
     end
    always @(m_mac_src_0_s0_27)
     begin
      mac_src_0_s0_27 <= m_mac_src_0_s0_27;
     end
    always @(m_mac_src_0_s0_28)
     begin
      mac_src_0_s0_28 <= m_mac_src_0_s0_28;
     end
    always @(m_mac_src_0_s0_29)
     begin
      mac_src_0_s0_29 <= m_mac_src_0_s0_29;
     end
    always @(m_mac_src_0_s0_30)
     begin
      mac_src_0_s0_30 <= m_mac_src_0_s0_30;
     end
    always @(m_mac_src_0_s0_31)
     begin
      mac_src_0_s0_31 <= m_mac_src_0_s0_31;
     end
    always @(m_mac_src_0_s1_0)
     begin
      mac_src_0_s1_0 <= m_mac_src_0_s1_0;
     end
    always @(m_mac_src_0_s1_1)
     begin
      mac_src_0_s1_1 <= m_mac_src_0_s1_1;
     end
    always @(m_mac_src_0_s1_2)
     begin
      mac_src_0_s1_2 <= m_mac_src_0_s1_2;
     end
    always @(m_mac_src_0_s1_3)
     begin
      mac_src_0_s1_3 <= m_mac_src_0_s1_3;
     end
    always @(m_mac_src_0_s1_4)
     begin
      mac_src_0_s1_4 <= m_mac_src_0_s1_4;
     end
    always @(m_mac_src_0_s1_5)
     begin
      mac_src_0_s1_5 <= m_mac_src_0_s1_5;
     end
    always @(m_mac_src_0_s1_6)
     begin
      mac_src_0_s1_6 <= m_mac_src_0_s1_6;
     end
    always @(m_mac_src_0_s1_7)
     begin
      mac_src_0_s1_7 <= m_mac_src_0_s1_7;
     end
    always @(m_mac_src_0_s1_8)
     begin
      mac_src_0_s1_8 <= m_mac_src_0_s1_8;
     end
    always @(m_mac_src_0_s1_9)
     begin
      mac_src_0_s1_9 <= m_mac_src_0_s1_9;
     end
    always @(m_mac_src_0_s1_10)
     begin
      mac_src_0_s1_10 <= m_mac_src_0_s1_10;
     end
    always @(m_mac_src_0_s1_11)
     begin
      mac_src_0_s1_11 <= m_mac_src_0_s1_11;
     end
    always @(m_mac_src_0_s1_12)
     begin
      mac_src_0_s1_12 <= m_mac_src_0_s1_12;
     end
    always @(m_mac_src_0_s1_13)
     begin
      mac_src_0_s1_13 <= m_mac_src_0_s1_13;
     end
    always @(m_mac_src_0_s1_14)
     begin
      mac_src_0_s1_14 <= m_mac_src_0_s1_14;
     end
    always @(m_mac_src_0_s1_15)
     begin
      mac_src_0_s1_15 <= m_mac_src_0_s1_15;
     end
    always @(m_mac_src_0_s1_16)
     begin
      mac_src_0_s1_16 <= m_mac_src_0_s1_16;
     end
    always @(m_mac_src_0_s1_17)
     begin
      mac_src_0_s1_17 <= m_mac_src_0_s1_17;
     end
    always @(m_mac_src_0_s1_18)
     begin
      mac_src_0_s1_18 <= m_mac_src_0_s1_18;
     end
    always @(m_mac_src_0_s1_19)
     begin
      mac_src_0_s1_19 <= m_mac_src_0_s1_19;
     end
    always @(m_mac_src_0_s1_20)
     begin
      mac_src_0_s1_20 <= m_mac_src_0_s1_20;
     end
    always @(m_mac_src_0_s1_21)
     begin
      mac_src_0_s1_21 <= m_mac_src_0_s1_21;
     end
    always @(m_mac_src_0_s1_22)
     begin
      mac_src_0_s1_22 <= m_mac_src_0_s1_22;
     end
    always @(m_mac_src_0_s1_23)
     begin
      mac_src_0_s1_23 <= m_mac_src_0_s1_23;
     end
    always @(m_mac_src_0_s1_24)
     begin
      mac_src_0_s1_24 <= m_mac_src_0_s1_24;
     end
    always @(m_mac_src_0_s1_25)
     begin
      mac_src_0_s1_25 <= m_mac_src_0_s1_25;
     end
    always @(m_mac_src_0_s1_26)
     begin
      mac_src_0_s1_26 <= m_mac_src_0_s1_26;
     end
    always @(m_mac_src_0_s1_27)
     begin
      mac_src_0_s1_27 <= m_mac_src_0_s1_27;
     end
    always @(m_mac_src_0_s1_28)
     begin
      mac_src_0_s1_28 <= m_mac_src_0_s1_28;
     end
    always @(m_mac_src_0_s1_29)
     begin
      mac_src_0_s1_29 <= m_mac_src_0_s1_29;
     end
    always @(m_mac_src_0_s1_30)
     begin
      mac_src_0_s1_30 <= m_mac_src_0_s1_30;
     end
    always @(m_mac_src_0_s1_31)
     begin
      mac_src_0_s1_31 <= m_mac_src_0_s1_31;
     end
    always @(m_mac_src_0_s2_0)
     begin
      mac_src_0_s2_0 <= m_mac_src_0_s2_0;
     end
    always @(m_mac_src_0_s2_1)
     begin
      mac_src_0_s2_1 <= m_mac_src_0_s2_1;
     end
    always @(m_mac_src_0_s2_2)
     begin
      mac_src_0_s2_2 <= m_mac_src_0_s2_2;
     end
    always @(m_mac_src_0_s2_3)
     begin
      mac_src_0_s2_3 <= m_mac_src_0_s2_3;
     end
    always @(m_mac_src_0_s2_4)
     begin
      mac_src_0_s2_4 <= m_mac_src_0_s2_4;
     end
    always @(m_mac_src_0_s2_5)
     begin
      mac_src_0_s2_5 <= m_mac_src_0_s2_5;
     end
    always @(m_mac_src_0_s2_6)
     begin
      mac_src_0_s2_6 <= m_mac_src_0_s2_6;
     end
    always @(m_mac_src_0_s2_7)
     begin
      mac_src_0_s2_7 <= m_mac_src_0_s2_7;
     end
    always @(m_mac_src_0_s2_8)
     begin
      mac_src_0_s2_8 <= m_mac_src_0_s2_8;
     end
    always @(m_mac_src_0_s2_9)
     begin
      mac_src_0_s2_9 <= m_mac_src_0_s2_9;
     end
    always @(m_mac_src_0_s2_10)
     begin
      mac_src_0_s2_10 <= m_mac_src_0_s2_10;
     end
    always @(m_mac_src_0_s2_11)
     begin
      mac_src_0_s2_11 <= m_mac_src_0_s2_11;
     end
    always @(m_mac_src_0_s2_12)
     begin
      mac_src_0_s2_12 <= m_mac_src_0_s2_12;
     end
    always @(m_mac_src_0_s2_13)
     begin
      mac_src_0_s2_13 <= m_mac_src_0_s2_13;
     end
    always @(m_mac_src_0_s2_14)
     begin
      mac_src_0_s2_14 <= m_mac_src_0_s2_14;
     end
    always @(m_mac_src_0_s2_15)
     begin
      mac_src_0_s2_15 <= m_mac_src_0_s2_15;
     end
    always @(m_mac_src_0_s2_16)
     begin
      mac_src_0_s2_16 <= m_mac_src_0_s2_16;
     end
    always @(m_mac_src_0_s2_17)
     begin
      mac_src_0_s2_17 <= m_mac_src_0_s2_17;
     end
    always @(m_mac_src_0_s2_18)
     begin
      mac_src_0_s2_18 <= m_mac_src_0_s2_18;
     end
    always @(m_mac_src_0_s2_19)
     begin
      mac_src_0_s2_19 <= m_mac_src_0_s2_19;
     end
    always @(m_mac_src_0_s2_20)
     begin
      mac_src_0_s2_20 <= m_mac_src_0_s2_20;
     end
    always @(m_mac_src_0_s2_21)
     begin
      mac_src_0_s2_21 <= m_mac_src_0_s2_21;
     end
    always @(m_mac_src_0_s2_22)
     begin
      mac_src_0_s2_22 <= m_mac_src_0_s2_22;
     end
    always @(m_mac_src_0_s2_23)
     begin
      mac_src_0_s2_23 <= m_mac_src_0_s2_23;
     end
    always @(m_mac_src_0_s2_24)
     begin
      mac_src_0_s2_24 <= m_mac_src_0_s2_24;
     end
    always @(m_mac_src_0_s2_25)
     begin
      mac_src_0_s2_25 <= m_mac_src_0_s2_25;
     end
    always @(m_mac_src_0_s2_26)
     begin
      mac_src_0_s2_26 <= m_mac_src_0_s2_26;
     end
    always @(m_mac_src_0_s2_27)
     begin
      mac_src_0_s2_27 <= m_mac_src_0_s2_27;
     end
    always @(m_mac_src_0_s2_28)
     begin
      mac_src_0_s2_28 <= m_mac_src_0_s2_28;
     end
    always @(m_mac_src_0_s2_29)
     begin
      mac_src_0_s2_29 <= m_mac_src_0_s2_29;
     end
    always @(m_mac_src_0_s2_30)
     begin
      mac_src_0_s2_30 <= m_mac_src_0_s2_30;
     end
    always @(m_mac_src_0_s2_31)
     begin
      mac_src_0_s2_31 <= m_mac_src_0_s2_31;
     end
    always @(m_mac_src_0_s3_0)
     begin
      mac_src_0_s3_0 <= m_mac_src_0_s3_0;
     end
    always @(m_mac_src_0_s3_1)
     begin
      mac_src_0_s3_1 <= m_mac_src_0_s3_1;
     end
    always @(m_mac_src_0_s3_2)
     begin
      mac_src_0_s3_2 <= m_mac_src_0_s3_2;
     end
    always @(m_mac_src_0_s3_3)
     begin
      mac_src_0_s3_3 <= m_mac_src_0_s3_3;
     end
    always @(m_mac_src_0_s3_4)
     begin
      mac_src_0_s3_4 <= m_mac_src_0_s3_4;
     end
    always @(m_mac_src_0_s3_5)
     begin
      mac_src_0_s3_5 <= m_mac_src_0_s3_5;
     end
    always @(m_mac_src_0_s3_6)
     begin
      mac_src_0_s3_6 <= m_mac_src_0_s3_6;
     end
    always @(m_mac_src_0_s3_7)
     begin
      mac_src_0_s3_7 <= m_mac_src_0_s3_7;
     end
    always @(m_mac_src_0_s3_8)
     begin
      mac_src_0_s3_8 <= m_mac_src_0_s3_8;
     end
    always @(m_mac_src_0_s3_9)
     begin
      mac_src_0_s3_9 <= m_mac_src_0_s3_9;
     end
    always @(m_mac_src_0_s3_10)
     begin
      mac_src_0_s3_10 <= m_mac_src_0_s3_10;
     end
    always @(m_mac_src_0_s3_11)
     begin
      mac_src_0_s3_11 <= m_mac_src_0_s3_11;
     end
    always @(m_mac_src_0_s3_12)
     begin
      mac_src_0_s3_12 <= m_mac_src_0_s3_12;
     end
    always @(m_mac_src_0_s3_13)
     begin
      mac_src_0_s3_13 <= m_mac_src_0_s3_13;
     end
    always @(m_mac_src_0_s3_14)
     begin
      mac_src_0_s3_14 <= m_mac_src_0_s3_14;
     end
    always @(m_mac_src_0_s3_15)
     begin
      mac_src_0_s3_15 <= m_mac_src_0_s3_15;
     end
    always @(m_mac_src_0_s3_16)
     begin
      mac_src_0_s3_16 <= m_mac_src_0_s3_16;
     end
    always @(m_mac_src_0_s3_17)
     begin
      mac_src_0_s3_17 <= m_mac_src_0_s3_17;
     end
    always @(m_mac_src_0_s3_18)
     begin
      mac_src_0_s3_18 <= m_mac_src_0_s3_18;
     end
    always @(m_mac_src_0_s3_19)
     begin
      mac_src_0_s3_19 <= m_mac_src_0_s3_19;
     end
    always @(m_mac_src_0_s3_20)
     begin
      mac_src_0_s3_20 <= m_mac_src_0_s3_20;
     end
    always @(m_mac_src_0_s3_21)
     begin
      mac_src_0_s3_21 <= m_mac_src_0_s3_21;
     end
    always @(m_mac_src_0_s3_22)
     begin
      mac_src_0_s3_22 <= m_mac_src_0_s3_22;
     end
    always @(m_mac_src_0_s3_23)
     begin
      mac_src_0_s3_23 <= m_mac_src_0_s3_23;
     end
    always @(m_mac_src_0_s3_24)
     begin
      mac_src_0_s3_24 <= m_mac_src_0_s3_24;
     end
    always @(m_mac_src_0_s3_25)
     begin
      mac_src_0_s3_25 <= m_mac_src_0_s3_25;
     end
    always @(m_mac_src_0_s3_26)
     begin
      mac_src_0_s3_26 <= m_mac_src_0_s3_26;
     end
    always @(m_mac_src_0_s3_27)
     begin
      mac_src_0_s3_27 <= m_mac_src_0_s3_27;
     end
    always @(m_mac_src_0_s3_28)
     begin
      mac_src_0_s3_28 <= m_mac_src_0_s3_28;
     end
    always @(m_mac_src_0_s3_29)
     begin
      mac_src_0_s3_29 <= m_mac_src_0_s3_29;
     end
    always @(m_mac_src_0_s3_30)
     begin
      mac_src_0_s3_30 <= m_mac_src_0_s3_30;
     end
    always @(m_mac_src_0_s3_31)
     begin
      mac_src_0_s3_31 <= m_mac_src_0_s3_31;
     end
    always @(m_mac_src_0_s4_0)
     begin
      mac_src_0_s4_0 <= m_mac_src_0_s4_0;
     end
    always @(m_mac_src_0_s4_1)
     begin
      mac_src_0_s4_1 <= m_mac_src_0_s4_1;
     end
    always @(m_mac_src_0_s4_2)
     begin
      mac_src_0_s4_2 <= m_mac_src_0_s4_2;
     end
    always @(m_mac_src_0_s4_3)
     begin
      mac_src_0_s4_3 <= m_mac_src_0_s4_3;
     end
    always @(m_mac_src_0_s4_4)
     begin
      mac_src_0_s4_4 <= m_mac_src_0_s4_4;
     end
    always @(m_mac_src_0_s4_5)
     begin
      mac_src_0_s4_5 <= m_mac_src_0_s4_5;
     end
    always @(m_mac_src_0_s4_6)
     begin
      mac_src_0_s4_6 <= m_mac_src_0_s4_6;
     end
    always @(m_mac_src_0_s4_7)
     begin
      mac_src_0_s4_7 <= m_mac_src_0_s4_7;
     end
    always @(m_mac_src_0_s4_8)
     begin
      mac_src_0_s4_8 <= m_mac_src_0_s4_8;
     end
    always @(m_mac_src_0_s4_9)
     begin
      mac_src_0_s4_9 <= m_mac_src_0_s4_9;
     end
    always @(m_mac_src_0_s4_10)
     begin
      mac_src_0_s4_10 <= m_mac_src_0_s4_10;
     end
    always @(m_mac_src_0_s4_11)
     begin
      mac_src_0_s4_11 <= m_mac_src_0_s4_11;
     end
    always @(m_mac_src_0_s4_12)
     begin
      mac_src_0_s4_12 <= m_mac_src_0_s4_12;
     end
    always @(m_mac_src_0_s4_13)
     begin
      mac_src_0_s4_13 <= m_mac_src_0_s4_13;
     end
    always @(m_mac_src_0_s4_14)
     begin
      mac_src_0_s4_14 <= m_mac_src_0_s4_14;
     end
    always @(m_mac_src_0_s4_15)
     begin
      mac_src_0_s4_15 <= m_mac_src_0_s4_15;
     end
    always @(m_mac_src_0_s4_16)
     begin
      mac_src_0_s4_16 <= m_mac_src_0_s4_16;
     end
    always @(m_mac_src_0_s4_17)
     begin
      mac_src_0_s4_17 <= m_mac_src_0_s4_17;
     end
    always @(m_mac_src_0_s4_18)
     begin
      mac_src_0_s4_18 <= m_mac_src_0_s4_18;
     end
    always @(m_mac_src_0_s4_19)
     begin
      mac_src_0_s4_19 <= m_mac_src_0_s4_19;
     end
    always @(m_mac_src_0_s4_20)
     begin
      mac_src_0_s4_20 <= m_mac_src_0_s4_20;
     end
    always @(m_mac_src_0_s4_21)
     begin
      mac_src_0_s4_21 <= m_mac_src_0_s4_21;
     end
    always @(m_mac_src_0_s4_22)
     begin
      mac_src_0_s4_22 <= m_mac_src_0_s4_22;
     end
    always @(m_mac_src_0_s4_23)
     begin
      mac_src_0_s4_23 <= m_mac_src_0_s4_23;
     end
    always @(m_mac_src_0_s4_24)
     begin
      mac_src_0_s4_24 <= m_mac_src_0_s4_24;
     end
    always @(m_mac_src_0_s4_25)
     begin
      mac_src_0_s4_25 <= m_mac_src_0_s4_25;
     end
    always @(m_mac_src_0_s4_26)
     begin
      mac_src_0_s4_26 <= m_mac_src_0_s4_26;
     end
    always @(m_mac_src_0_s4_27)
     begin
      mac_src_0_s4_27 <= m_mac_src_0_s4_27;
     end
    always @(m_mac_src_0_s4_28)
     begin
      mac_src_0_s4_28 <= m_mac_src_0_s4_28;
     end
    always @(m_mac_src_0_s4_29)
     begin
      mac_src_0_s4_29 <= m_mac_src_0_s4_29;
     end
    always @(m_mac_src_0_s4_30)
     begin
      mac_src_0_s4_30 <= m_mac_src_0_s4_30;
     end
    always @(m_mac_src_0_s4_31)
     begin
      mac_src_0_s4_31 <= m_mac_src_0_s4_31;
     end
    always @(m_mac_src_0_s5_0)
     begin
      mac_src_0_s5_0 <= m_mac_src_0_s5_0;
     end
    always @(m_mac_src_0_s5_1)
     begin
      mac_src_0_s5_1 <= m_mac_src_0_s5_1;
     end
    always @(m_mac_src_0_s5_2)
     begin
      mac_src_0_s5_2 <= m_mac_src_0_s5_2;
     end
    always @(m_mac_src_0_s5_3)
     begin
      mac_src_0_s5_3 <= m_mac_src_0_s5_3;
     end
    always @(m_mac_src_0_s5_4)
     begin
      mac_src_0_s5_4 <= m_mac_src_0_s5_4;
     end
    always @(m_mac_src_0_s5_5)
     begin
      mac_src_0_s5_5 <= m_mac_src_0_s5_5;
     end
    always @(m_mac_src_0_s5_6)
     begin
      mac_src_0_s5_6 <= m_mac_src_0_s5_6;
     end
    always @(m_mac_src_0_s5_7)
     begin
      mac_src_0_s5_7 <= m_mac_src_0_s5_7;
     end
    always @(m_mac_src_0_s5_8)
     begin
      mac_src_0_s5_8 <= m_mac_src_0_s5_8;
     end
    always @(m_mac_src_0_s5_9)
     begin
      mac_src_0_s5_9 <= m_mac_src_0_s5_9;
     end
    always @(m_mac_src_0_s5_10)
     begin
      mac_src_0_s5_10 <= m_mac_src_0_s5_10;
     end
    always @(m_mac_src_0_s5_11)
     begin
      mac_src_0_s5_11 <= m_mac_src_0_s5_11;
     end
    always @(m_mac_src_0_s5_12)
     begin
      mac_src_0_s5_12 <= m_mac_src_0_s5_12;
     end
    always @(m_mac_src_0_s5_13)
     begin
      mac_src_0_s5_13 <= m_mac_src_0_s5_13;
     end
    always @(m_mac_src_0_s5_14)
     begin
      mac_src_0_s5_14 <= m_mac_src_0_s5_14;
     end
    always @(m_mac_src_0_s5_15)
     begin
      mac_src_0_s5_15 <= m_mac_src_0_s5_15;
     end
    always @(m_mac_src_0_s5_16)
     begin
      mac_src_0_s5_16 <= m_mac_src_0_s5_16;
     end
    always @(m_mac_src_0_s5_17)
     begin
      mac_src_0_s5_17 <= m_mac_src_0_s5_17;
     end
    always @(m_mac_src_0_s5_18)
     begin
      mac_src_0_s5_18 <= m_mac_src_0_s5_18;
     end
    always @(m_mac_src_0_s5_19)
     begin
      mac_src_0_s5_19 <= m_mac_src_0_s5_19;
     end
    always @(m_mac_src_0_s5_20)
     begin
      mac_src_0_s5_20 <= m_mac_src_0_s5_20;
     end
    always @(m_mac_src_0_s5_21)
     begin
      mac_src_0_s5_21 <= m_mac_src_0_s5_21;
     end
    always @(m_mac_src_0_s5_22)
     begin
      mac_src_0_s5_22 <= m_mac_src_0_s5_22;
     end
    always @(m_mac_src_0_s5_23)
     begin
      mac_src_0_s5_23 <= m_mac_src_0_s5_23;
     end
    always @(m_mac_src_0_s5_24)
     begin
      mac_src_0_s5_24 <= m_mac_src_0_s5_24;
     end
    always @(m_mac_src_0_s5_25)
     begin
      mac_src_0_s5_25 <= m_mac_src_0_s5_25;
     end
    always @(m_mac_src_0_s5_26)
     begin
      mac_src_0_s5_26 <= m_mac_src_0_s5_26;
     end
    always @(m_mac_src_0_s5_27)
     begin
      mac_src_0_s5_27 <= m_mac_src_0_s5_27;
     end
    always @(m_mac_src_0_s5_28)
     begin
      mac_src_0_s5_28 <= m_mac_src_0_s5_28;
     end
    always @(m_mac_src_0_s5_29)
     begin
      mac_src_0_s5_29 <= m_mac_src_0_s5_29;
     end
    always @(m_mac_src_0_s5_30)
     begin
      mac_src_0_s5_30 <= m_mac_src_0_s5_30;
     end
    always @(m_mac_src_0_s5_31)
     begin
      mac_src_0_s5_31 <= m_mac_src_0_s5_31;
     end
    always @(m_mac_src_0_s6_0)
     begin
      mac_src_0_s6_0 <= m_mac_src_0_s6_0;
     end
    always @(m_mac_src_0_s6_1)
     begin
      mac_src_0_s6_1 <= m_mac_src_0_s6_1;
     end
    always @(m_mac_src_0_s6_2)
     begin
      mac_src_0_s6_2 <= m_mac_src_0_s6_2;
     end
    always @(m_mac_src_0_s6_3)
     begin
      mac_src_0_s6_3 <= m_mac_src_0_s6_3;
     end
    always @(m_mac_src_0_s6_4)
     begin
      mac_src_0_s6_4 <= m_mac_src_0_s6_4;
     end
    always @(m_mac_src_0_s6_5)
     begin
      mac_src_0_s6_5 <= m_mac_src_0_s6_5;
     end
    always @(m_mac_src_0_s6_6)
     begin
      mac_src_0_s6_6 <= m_mac_src_0_s6_6;
     end
    always @(m_mac_src_0_s6_7)
     begin
      mac_src_0_s6_7 <= m_mac_src_0_s6_7;
     end
    always @(m_mac_src_0_s6_8)
     begin
      mac_src_0_s6_8 <= m_mac_src_0_s6_8;
     end
    always @(m_mac_src_0_s6_9)
     begin
      mac_src_0_s6_9 <= m_mac_src_0_s6_9;
     end
    always @(m_mac_src_0_s6_10)
     begin
      mac_src_0_s6_10 <= m_mac_src_0_s6_10;
     end
    always @(m_mac_src_0_s6_11)
     begin
      mac_src_0_s6_11 <= m_mac_src_0_s6_11;
     end
    always @(m_mac_src_0_s6_12)
     begin
      mac_src_0_s6_12 <= m_mac_src_0_s6_12;
     end
    always @(m_mac_src_0_s6_13)
     begin
      mac_src_0_s6_13 <= m_mac_src_0_s6_13;
     end
    always @(m_mac_src_0_s6_14)
     begin
      mac_src_0_s6_14 <= m_mac_src_0_s6_14;
     end
    always @(m_mac_src_0_s6_15)
     begin
      mac_src_0_s6_15 <= m_mac_src_0_s6_15;
     end
    always @(m_mac_src_0_s6_16)
     begin
      mac_src_0_s6_16 <= m_mac_src_0_s6_16;
     end
    always @(m_mac_src_0_s6_17)
     begin
      mac_src_0_s6_17 <= m_mac_src_0_s6_17;
     end
    always @(m_mac_src_0_s6_18)
     begin
      mac_src_0_s6_18 <= m_mac_src_0_s6_18;
     end
    always @(m_mac_src_0_s6_19)
     begin
      mac_src_0_s6_19 <= m_mac_src_0_s6_19;
     end
    always @(m_mac_src_0_s6_20)
     begin
      mac_src_0_s6_20 <= m_mac_src_0_s6_20;
     end
    always @(m_mac_src_0_s6_21)
     begin
      mac_src_0_s6_21 <= m_mac_src_0_s6_21;
     end
    always @(m_mac_src_0_s6_22)
     begin
      mac_src_0_s6_22 <= m_mac_src_0_s6_22;
     end
    always @(m_mac_src_0_s6_23)
     begin
      mac_src_0_s6_23 <= m_mac_src_0_s6_23;
     end
    always @(m_mac_src_0_s6_24)
     begin
      mac_src_0_s6_24 <= m_mac_src_0_s6_24;
     end
    always @(m_mac_src_0_s6_25)
     begin
      mac_src_0_s6_25 <= m_mac_src_0_s6_25;
     end
    always @(m_mac_src_0_s6_26)
     begin
      mac_src_0_s6_26 <= m_mac_src_0_s6_26;
     end
    always @(m_mac_src_0_s6_27)
     begin
      mac_src_0_s6_27 <= m_mac_src_0_s6_27;
     end
    always @(m_mac_src_0_s6_28)
     begin
      mac_src_0_s6_28 <= m_mac_src_0_s6_28;
     end
    always @(m_mac_src_0_s6_29)
     begin
      mac_src_0_s6_29 <= m_mac_src_0_s6_29;
     end
    always @(m_mac_src_0_s6_30)
     begin
      mac_src_0_s6_30 <= m_mac_src_0_s6_30;
     end
    always @(m_mac_src_0_s6_31)
     begin
      mac_src_0_s6_31 <= m_mac_src_0_s6_31;
     end
    always @(m_mac_src_1_0)
     begin
      mac_src_1_0 <= m_mac_src_1_0;
     end
    always @(m_mac_src_1_1)
     begin
      mac_src_1_1 <= m_mac_src_1_1;
     end
    always @(m_mac_src_1_2)
     begin
      mac_src_1_2 <= m_mac_src_1_2;
     end
    always @(m_mac_src_1_3)
     begin
      mac_src_1_3 <= m_mac_src_1_3;
     end
    always @(m_mac_src_1_4)
     begin
      mac_src_1_4 <= m_mac_src_1_4;
     end
    always @(m_mac_src_1_5)
     begin
      mac_src_1_5 <= m_mac_src_1_5;
     end
    always @(m_mac_src_1_6)
     begin
      mac_src_1_6 <= m_mac_src_1_6;
     end
    always @(m_mac_src_1_7)
     begin
      mac_src_1_7 <= m_mac_src_1_7;
     end
    always @(m_mac_src_1_8)
     begin
      mac_src_1_8 <= m_mac_src_1_8;
     end
    always @(m_mac_src_1_9)
     begin
      mac_src_1_9 <= m_mac_src_1_9;
     end
    always @(m_mac_src_1_10)
     begin
      mac_src_1_10 <= m_mac_src_1_10;
     end
    always @(m_mac_src_1_11)
     begin
      mac_src_1_11 <= m_mac_src_1_11;
     end
    always @(m_mac_src_1_12)
     begin
      mac_src_1_12 <= m_mac_src_1_12;
     end
    always @(m_mac_src_1_13)
     begin
      mac_src_1_13 <= m_mac_src_1_13;
     end
    always @(m_mac_src_1_14)
     begin
      mac_src_1_14 <= m_mac_src_1_14;
     end
    always @(m_mac_src_1_15)
     begin
      mac_src_1_15 <= m_mac_src_1_15;
     end
    always @(m_mac_src_1_16)
     begin
      mac_src_1_16 <= m_mac_src_1_16;
     end
    always @(m_mac_src_1_17)
     begin
      mac_src_1_17 <= m_mac_src_1_17;
     end
    always @(m_mac_src_1_18)
     begin
      mac_src_1_18 <= m_mac_src_1_18;
     end
    always @(m_mac_src_1_19)
     begin
      mac_src_1_19 <= m_mac_src_1_19;
     end
    always @(m_mac_src_1_20)
     begin
      mac_src_1_20 <= m_mac_src_1_20;
     end
    always @(m_mac_src_1_21)
     begin
      mac_src_1_21 <= m_mac_src_1_21;
     end
    always @(m_mac_src_1_22)
     begin
      mac_src_1_22 <= m_mac_src_1_22;
     end
    always @(m_mac_src_1_23)
     begin
      mac_src_1_23 <= m_mac_src_1_23;
     end
    always @(m_mac_src_1_24)
     begin
      mac_src_1_24 <= m_mac_src_1_24;
     end
    always @(m_mac_src_1_25)
     begin
      mac_src_1_25 <= m_mac_src_1_25;
     end
    always @(m_mac_src_1_26)
     begin
      mac_src_1_26 <= m_mac_src_1_26;
     end
    always @(m_mac_src_1_27)
     begin
      mac_src_1_27 <= m_mac_src_1_27;
     end
    always @(m_mac_src_1_28)
     begin
      mac_src_1_28 <= m_mac_src_1_28;
     end
    always @(m_mac_src_1_29)
     begin
      mac_src_1_29 <= m_mac_src_1_29;
     end
    always @(m_mac_src_1_30)
     begin
      mac_src_1_30 <= m_mac_src_1_30;
     end
    always @(m_mac_src_1_31)
     begin
      mac_src_1_31 <= m_mac_src_1_31;
     end
    always @(m_mac_src_valid)
     begin
      mac_src_valid <= m_mac_src_valid;
     end
    always @(m_mac_clear)
     begin
      mac_clear <= m_mac_clear;
     end


endmodule

// This is an internal module that instantiates the user's SystemC input module
// using the Incisive foreign module instantiation feature.
// The name of the module and the names of the inputs and outputs must match
// with those defined in the SystemC type_wrapper module
module cache_type_wrapper(
      clk,
       rstn,
       cache_en,
       systolic_en,
       systolic_depth,
       addr_if_start,
       systolic_sel,
       feature_data,
       feature_share_en,
       feature_data_en,
       feature_data_sel,
       weight_data,
       weight_data_en,
       mac_src_0_s0_0,
      mac_src_0_s0_1,
      mac_src_0_s0_2,
      mac_src_0_s0_3,
      mac_src_0_s0_4,
      mac_src_0_s0_5,
      mac_src_0_s0_6,
      mac_src_0_s0_7,
      mac_src_0_s0_8,
      mac_src_0_s0_9,
      mac_src_0_s0_10,
      mac_src_0_s0_11,
      mac_src_0_s0_12,
      mac_src_0_s0_13,
      mac_src_0_s0_14,
      mac_src_0_s0_15,
      mac_src_0_s0_16,
      mac_src_0_s0_17,
      mac_src_0_s0_18,
      mac_src_0_s0_19,
      mac_src_0_s0_20,
      mac_src_0_s0_21,
      mac_src_0_s0_22,
      mac_src_0_s0_23,
      mac_src_0_s0_24,
      mac_src_0_s0_25,
      mac_src_0_s0_26,
      mac_src_0_s0_27,
      mac_src_0_s0_28,
      mac_src_0_s0_29,
      mac_src_0_s0_30,
      mac_src_0_s0_31,
       mac_src_0_s1_0,
      mac_src_0_s1_1,
      mac_src_0_s1_2,
      mac_src_0_s1_3,
      mac_src_0_s1_4,
      mac_src_0_s1_5,
      mac_src_0_s1_6,
      mac_src_0_s1_7,
      mac_src_0_s1_8,
      mac_src_0_s1_9,
      mac_src_0_s1_10,
      mac_src_0_s1_11,
      mac_src_0_s1_12,
      mac_src_0_s1_13,
      mac_src_0_s1_14,
      mac_src_0_s1_15,
      mac_src_0_s1_16,
      mac_src_0_s1_17,
      mac_src_0_s1_18,
      mac_src_0_s1_19,
      mac_src_0_s1_20,
      mac_src_0_s1_21,
      mac_src_0_s1_22,
      mac_src_0_s1_23,
      mac_src_0_s1_24,
      mac_src_0_s1_25,
      mac_src_0_s1_26,
      mac_src_0_s1_27,
      mac_src_0_s1_28,
      mac_src_0_s1_29,
      mac_src_0_s1_30,
      mac_src_0_s1_31,
       mac_src_0_s2_0,
      mac_src_0_s2_1,
      mac_src_0_s2_2,
      mac_src_0_s2_3,
      mac_src_0_s2_4,
      mac_src_0_s2_5,
      mac_src_0_s2_6,
      mac_src_0_s2_7,
      mac_src_0_s2_8,
      mac_src_0_s2_9,
      mac_src_0_s2_10,
      mac_src_0_s2_11,
      mac_src_0_s2_12,
      mac_src_0_s2_13,
      mac_src_0_s2_14,
      mac_src_0_s2_15,
      mac_src_0_s2_16,
      mac_src_0_s2_17,
      mac_src_0_s2_18,
      mac_src_0_s2_19,
      mac_src_0_s2_20,
      mac_src_0_s2_21,
      mac_src_0_s2_22,
      mac_src_0_s2_23,
      mac_src_0_s2_24,
      mac_src_0_s2_25,
      mac_src_0_s2_26,
      mac_src_0_s2_27,
      mac_src_0_s2_28,
      mac_src_0_s2_29,
      mac_src_0_s2_30,
      mac_src_0_s2_31,
       mac_src_0_s3_0,
      mac_src_0_s3_1,
      mac_src_0_s3_2,
      mac_src_0_s3_3,
      mac_src_0_s3_4,
      mac_src_0_s3_5,
      mac_src_0_s3_6,
      mac_src_0_s3_7,
      mac_src_0_s3_8,
      mac_src_0_s3_9,
      mac_src_0_s3_10,
      mac_src_0_s3_11,
      mac_src_0_s3_12,
      mac_src_0_s3_13,
      mac_src_0_s3_14,
      mac_src_0_s3_15,
      mac_src_0_s3_16,
      mac_src_0_s3_17,
      mac_src_0_s3_18,
      mac_src_0_s3_19,
      mac_src_0_s3_20,
      mac_src_0_s3_21,
      mac_src_0_s3_22,
      mac_src_0_s3_23,
      mac_src_0_s3_24,
      mac_src_0_s3_25,
      mac_src_0_s3_26,
      mac_src_0_s3_27,
      mac_src_0_s3_28,
      mac_src_0_s3_29,
      mac_src_0_s3_30,
      mac_src_0_s3_31,
       mac_src_0_s4_0,
      mac_src_0_s4_1,
      mac_src_0_s4_2,
      mac_src_0_s4_3,
      mac_src_0_s4_4,
      mac_src_0_s4_5,
      mac_src_0_s4_6,
      mac_src_0_s4_7,
      mac_src_0_s4_8,
      mac_src_0_s4_9,
      mac_src_0_s4_10,
      mac_src_0_s4_11,
      mac_src_0_s4_12,
      mac_src_0_s4_13,
      mac_src_0_s4_14,
      mac_src_0_s4_15,
      mac_src_0_s4_16,
      mac_src_0_s4_17,
      mac_src_0_s4_18,
      mac_src_0_s4_19,
      mac_src_0_s4_20,
      mac_src_0_s4_21,
      mac_src_0_s4_22,
      mac_src_0_s4_23,
      mac_src_0_s4_24,
      mac_src_0_s4_25,
      mac_src_0_s4_26,
      mac_src_0_s4_27,
      mac_src_0_s4_28,
      mac_src_0_s4_29,
      mac_src_0_s4_30,
      mac_src_0_s4_31,
       mac_src_0_s5_0,
      mac_src_0_s5_1,
      mac_src_0_s5_2,
      mac_src_0_s5_3,
      mac_src_0_s5_4,
      mac_src_0_s5_5,
      mac_src_0_s5_6,
      mac_src_0_s5_7,
      mac_src_0_s5_8,
      mac_src_0_s5_9,
      mac_src_0_s5_10,
      mac_src_0_s5_11,
      mac_src_0_s5_12,
      mac_src_0_s5_13,
      mac_src_0_s5_14,
      mac_src_0_s5_15,
      mac_src_0_s5_16,
      mac_src_0_s5_17,
      mac_src_0_s5_18,
      mac_src_0_s5_19,
      mac_src_0_s5_20,
      mac_src_0_s5_21,
      mac_src_0_s5_22,
      mac_src_0_s5_23,
      mac_src_0_s5_24,
      mac_src_0_s5_25,
      mac_src_0_s5_26,
      mac_src_0_s5_27,
      mac_src_0_s5_28,
      mac_src_0_s5_29,
      mac_src_0_s5_30,
      mac_src_0_s5_31,
       mac_src_0_s6_0,
      mac_src_0_s6_1,
      mac_src_0_s6_2,
      mac_src_0_s6_3,
      mac_src_0_s6_4,
      mac_src_0_s6_5,
      mac_src_0_s6_6,
      mac_src_0_s6_7,
      mac_src_0_s6_8,
      mac_src_0_s6_9,
      mac_src_0_s6_10,
      mac_src_0_s6_11,
      mac_src_0_s6_12,
      mac_src_0_s6_13,
      mac_src_0_s6_14,
      mac_src_0_s6_15,
      mac_src_0_s6_16,
      mac_src_0_s6_17,
      mac_src_0_s6_18,
      mac_src_0_s6_19,
      mac_src_0_s6_20,
      mac_src_0_s6_21,
      mac_src_0_s6_22,
      mac_src_0_s6_23,
      mac_src_0_s6_24,
      mac_src_0_s6_25,
      mac_src_0_s6_26,
      mac_src_0_s6_27,
      mac_src_0_s6_28,
      mac_src_0_s6_29,
      mac_src_0_s6_30,
      mac_src_0_s6_31,
       mac_src_1_0,
      mac_src_1_1,
      mac_src_1_2,
      mac_src_1_3,
      mac_src_1_4,
      mac_src_1_5,
      mac_src_1_6,
      mac_src_1_7,
      mac_src_1_8,
      mac_src_1_9,
      mac_src_1_10,
      mac_src_1_11,
      mac_src_1_12,
      mac_src_1_13,
      mac_src_1_14,
      mac_src_1_15,
      mac_src_1_16,
      mac_src_1_17,
      mac_src_1_18,
      mac_src_1_19,
      mac_src_1_20,
      mac_src_1_21,
      mac_src_1_22,
      mac_src_1_23,
      mac_src_1_24,
      mac_src_1_25,
      mac_src_1_26,
      mac_src_1_27,
      mac_src_1_28,
      mac_src_1_29,
      mac_src_1_30,
      mac_src_1_31,
       mac_src_valid,
       mac_clear

    ) (* integer foreign = "SystemC";
    *);

	input clk;
	input rstn;
	input cache_en;
	input [7:0] systolic_en;
	input [7:0] systolic_depth;
	input addr_if_start;
	input [7:0] systolic_sel;
	input [319:0] feature_data;
	input feature_share_en;
	input feature_data_en;
	input [15:0] feature_data_sel;
	input [255:0] weight_data;
	input weight_data_en;
	output [9:0] mac_src_0_s0_0;
	output [9:0] mac_src_0_s0_1;
	output [9:0] mac_src_0_s0_2;
	output [9:0] mac_src_0_s0_3;
	output [9:0] mac_src_0_s0_4;
	output [9:0] mac_src_0_s0_5;
	output [9:0] mac_src_0_s0_6;
	output [9:0] mac_src_0_s0_7;
	output [9:0] mac_src_0_s0_8;
	output [9:0] mac_src_0_s0_9;
	output [9:0] mac_src_0_s0_10;
	output [9:0] mac_src_0_s0_11;
	output [9:0] mac_src_0_s0_12;
	output [9:0] mac_src_0_s0_13;
	output [9:0] mac_src_0_s0_14;
	output [9:0] mac_src_0_s0_15;
	output [9:0] mac_src_0_s0_16;
	output [9:0] mac_src_0_s0_17;
	output [9:0] mac_src_0_s0_18;
	output [9:0] mac_src_0_s0_19;
	output [9:0] mac_src_0_s0_20;
	output [9:0] mac_src_0_s0_21;
	output [9:0] mac_src_0_s0_22;
	output [9:0] mac_src_0_s0_23;
	output [9:0] mac_src_0_s0_24;
	output [9:0] mac_src_0_s0_25;
	output [9:0] mac_src_0_s0_26;
	output [9:0] mac_src_0_s0_27;
	output [9:0] mac_src_0_s0_28;
	output [9:0] mac_src_0_s0_29;
	output [9:0] mac_src_0_s0_30;
	output [9:0] mac_src_0_s0_31;
	output [9:0] mac_src_0_s1_0;
	output [9:0] mac_src_0_s1_1;
	output [9:0] mac_src_0_s1_2;
	output [9:0] mac_src_0_s1_3;
	output [9:0] mac_src_0_s1_4;
	output [9:0] mac_src_0_s1_5;
	output [9:0] mac_src_0_s1_6;
	output [9:0] mac_src_0_s1_7;
	output [9:0] mac_src_0_s1_8;
	output [9:0] mac_src_0_s1_9;
	output [9:0] mac_src_0_s1_10;
	output [9:0] mac_src_0_s1_11;
	output [9:0] mac_src_0_s1_12;
	output [9:0] mac_src_0_s1_13;
	output [9:0] mac_src_0_s1_14;
	output [9:0] mac_src_0_s1_15;
	output [9:0] mac_src_0_s1_16;
	output [9:0] mac_src_0_s1_17;
	output [9:0] mac_src_0_s1_18;
	output [9:0] mac_src_0_s1_19;
	output [9:0] mac_src_0_s1_20;
	output [9:0] mac_src_0_s1_21;
	output [9:0] mac_src_0_s1_22;
	output [9:0] mac_src_0_s1_23;
	output [9:0] mac_src_0_s1_24;
	output [9:0] mac_src_0_s1_25;
	output [9:0] mac_src_0_s1_26;
	output [9:0] mac_src_0_s1_27;
	output [9:0] mac_src_0_s1_28;
	output [9:0] mac_src_0_s1_29;
	output [9:0] mac_src_0_s1_30;
	output [9:0] mac_src_0_s1_31;
	output [9:0] mac_src_0_s2_0;
	output [9:0] mac_src_0_s2_1;
	output [9:0] mac_src_0_s2_2;
	output [9:0] mac_src_0_s2_3;
	output [9:0] mac_src_0_s2_4;
	output [9:0] mac_src_0_s2_5;
	output [9:0] mac_src_0_s2_6;
	output [9:0] mac_src_0_s2_7;
	output [9:0] mac_src_0_s2_8;
	output [9:0] mac_src_0_s2_9;
	output [9:0] mac_src_0_s2_10;
	output [9:0] mac_src_0_s2_11;
	output [9:0] mac_src_0_s2_12;
	output [9:0] mac_src_0_s2_13;
	output [9:0] mac_src_0_s2_14;
	output [9:0] mac_src_0_s2_15;
	output [9:0] mac_src_0_s2_16;
	output [9:0] mac_src_0_s2_17;
	output [9:0] mac_src_0_s2_18;
	output [9:0] mac_src_0_s2_19;
	output [9:0] mac_src_0_s2_20;
	output [9:0] mac_src_0_s2_21;
	output [9:0] mac_src_0_s2_22;
	output [9:0] mac_src_0_s2_23;
	output [9:0] mac_src_0_s2_24;
	output [9:0] mac_src_0_s2_25;
	output [9:0] mac_src_0_s2_26;
	output [9:0] mac_src_0_s2_27;
	output [9:0] mac_src_0_s2_28;
	output [9:0] mac_src_0_s2_29;
	output [9:0] mac_src_0_s2_30;
	output [9:0] mac_src_0_s2_31;
	output [9:0] mac_src_0_s3_0;
	output [9:0] mac_src_0_s3_1;
	output [9:0] mac_src_0_s3_2;
	output [9:0] mac_src_0_s3_3;
	output [9:0] mac_src_0_s3_4;
	output [9:0] mac_src_0_s3_5;
	output [9:0] mac_src_0_s3_6;
	output [9:0] mac_src_0_s3_7;
	output [9:0] mac_src_0_s3_8;
	output [9:0] mac_src_0_s3_9;
	output [9:0] mac_src_0_s3_10;
	output [9:0] mac_src_0_s3_11;
	output [9:0] mac_src_0_s3_12;
	output [9:0] mac_src_0_s3_13;
	output [9:0] mac_src_0_s3_14;
	output [9:0] mac_src_0_s3_15;
	output [9:0] mac_src_0_s3_16;
	output [9:0] mac_src_0_s3_17;
	output [9:0] mac_src_0_s3_18;
	output [9:0] mac_src_0_s3_19;
	output [9:0] mac_src_0_s3_20;
	output [9:0] mac_src_0_s3_21;
	output [9:0] mac_src_0_s3_22;
	output [9:0] mac_src_0_s3_23;
	output [9:0] mac_src_0_s3_24;
	output [9:0] mac_src_0_s3_25;
	output [9:0] mac_src_0_s3_26;
	output [9:0] mac_src_0_s3_27;
	output [9:0] mac_src_0_s3_28;
	output [9:0] mac_src_0_s3_29;
	output [9:0] mac_src_0_s3_30;
	output [9:0] mac_src_0_s3_31;
	output [9:0] mac_src_0_s4_0;
	output [9:0] mac_src_0_s4_1;
	output [9:0] mac_src_0_s4_2;
	output [9:0] mac_src_0_s4_3;
	output [9:0] mac_src_0_s4_4;
	output [9:0] mac_src_0_s4_5;
	output [9:0] mac_src_0_s4_6;
	output [9:0] mac_src_0_s4_7;
	output [9:0] mac_src_0_s4_8;
	output [9:0] mac_src_0_s4_9;
	output [9:0] mac_src_0_s4_10;
	output [9:0] mac_src_0_s4_11;
	output [9:0] mac_src_0_s4_12;
	output [9:0] mac_src_0_s4_13;
	output [9:0] mac_src_0_s4_14;
	output [9:0] mac_src_0_s4_15;
	output [9:0] mac_src_0_s4_16;
	output [9:0] mac_src_0_s4_17;
	output [9:0] mac_src_0_s4_18;
	output [9:0] mac_src_0_s4_19;
	output [9:0] mac_src_0_s4_20;
	output [9:0] mac_src_0_s4_21;
	output [9:0] mac_src_0_s4_22;
	output [9:0] mac_src_0_s4_23;
	output [9:0] mac_src_0_s4_24;
	output [9:0] mac_src_0_s4_25;
	output [9:0] mac_src_0_s4_26;
	output [9:0] mac_src_0_s4_27;
	output [9:0] mac_src_0_s4_28;
	output [9:0] mac_src_0_s4_29;
	output [9:0] mac_src_0_s4_30;
	output [9:0] mac_src_0_s4_31;
	output [9:0] mac_src_0_s5_0;
	output [9:0] mac_src_0_s5_1;
	output [9:0] mac_src_0_s5_2;
	output [9:0] mac_src_0_s5_3;
	output [9:0] mac_src_0_s5_4;
	output [9:0] mac_src_0_s5_5;
	output [9:0] mac_src_0_s5_6;
	output [9:0] mac_src_0_s5_7;
	output [9:0] mac_src_0_s5_8;
	output [9:0] mac_src_0_s5_9;
	output [9:0] mac_src_0_s5_10;
	output [9:0] mac_src_0_s5_11;
	output [9:0] mac_src_0_s5_12;
	output [9:0] mac_src_0_s5_13;
	output [9:0] mac_src_0_s5_14;
	output [9:0] mac_src_0_s5_15;
	output [9:0] mac_src_0_s5_16;
	output [9:0] mac_src_0_s5_17;
	output [9:0] mac_src_0_s5_18;
	output [9:0] mac_src_0_s5_19;
	output [9:0] mac_src_0_s5_20;
	output [9:0] mac_src_0_s5_21;
	output [9:0] mac_src_0_s5_22;
	output [9:0] mac_src_0_s5_23;
	output [9:0] mac_src_0_s5_24;
	output [9:0] mac_src_0_s5_25;
	output [9:0] mac_src_0_s5_26;
	output [9:0] mac_src_0_s5_27;
	output [9:0] mac_src_0_s5_28;
	output [9:0] mac_src_0_s5_29;
	output [9:0] mac_src_0_s5_30;
	output [9:0] mac_src_0_s5_31;
	output [9:0] mac_src_0_s6_0;
	output [9:0] mac_src_0_s6_1;
	output [9:0] mac_src_0_s6_2;
	output [9:0] mac_src_0_s6_3;
	output [9:0] mac_src_0_s6_4;
	output [9:0] mac_src_0_s6_5;
	output [9:0] mac_src_0_s6_6;
	output [9:0] mac_src_0_s6_7;
	output [9:0] mac_src_0_s6_8;
	output [9:0] mac_src_0_s6_9;
	output [9:0] mac_src_0_s6_10;
	output [9:0] mac_src_0_s6_11;
	output [9:0] mac_src_0_s6_12;
	output [9:0] mac_src_0_s6_13;
	output [9:0] mac_src_0_s6_14;
	output [9:0] mac_src_0_s6_15;
	output [9:0] mac_src_0_s6_16;
	output [9:0] mac_src_0_s6_17;
	output [9:0] mac_src_0_s6_18;
	output [9:0] mac_src_0_s6_19;
	output [9:0] mac_src_0_s6_20;
	output [9:0] mac_src_0_s6_21;
	output [9:0] mac_src_0_s6_22;
	output [9:0] mac_src_0_s6_23;
	output [9:0] mac_src_0_s6_24;
	output [9:0] mac_src_0_s6_25;
	output [9:0] mac_src_0_s6_26;
	output [9:0] mac_src_0_s6_27;
	output [9:0] mac_src_0_s6_28;
	output [9:0] mac_src_0_s6_29;
	output [9:0] mac_src_0_s6_30;
	output [9:0] mac_src_0_s6_31;
	output [7:0] mac_src_1_0;
	output [7:0] mac_src_1_1;
	output [7:0] mac_src_1_2;
	output [7:0] mac_src_1_3;
	output [7:0] mac_src_1_4;
	output [7:0] mac_src_1_5;
	output [7:0] mac_src_1_6;
	output [7:0] mac_src_1_7;
	output [7:0] mac_src_1_8;
	output [7:0] mac_src_1_9;
	output [7:0] mac_src_1_10;
	output [7:0] mac_src_1_11;
	output [7:0] mac_src_1_12;
	output [7:0] mac_src_1_13;
	output [7:0] mac_src_1_14;
	output [7:0] mac_src_1_15;
	output [7:0] mac_src_1_16;
	output [7:0] mac_src_1_17;
	output [7:0] mac_src_1_18;
	output [7:0] mac_src_1_19;
	output [7:0] mac_src_1_20;
	output [7:0] mac_src_1_21;
	output [7:0] mac_src_1_22;
	output [7:0] mac_src_1_23;
	output [7:0] mac_src_1_24;
	output [7:0] mac_src_1_25;
	output [7:0] mac_src_1_26;
	output [7:0] mac_src_1_27;
	output [7:0] mac_src_1_28;
	output [7:0] mac_src_1_29;
	output [7:0] mac_src_1_30;
	output [7:0] mac_src_1_31;
	output mac_src_valid;
	output mac_clear;


endmodule
