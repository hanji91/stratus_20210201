/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:20 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2052368036_bdw (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__46,
	inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49,
	inst_cellmath__51;
wire N440,N441,N442,N443,N444,N445,N446 
	,N447,N448,N449,N450,N461,N462,N463,N469 
	,N470;
cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I0 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw2052368036_bdw cynw_cm_float_mul_ieee_I1 (.inst_cellmath__19__2__out0(inst_cellmath__19), .inst_cellmath__19__2__in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I2 (.inst_cellmath__21_0_out0(inst_cellmath__21), .inst_cellmath__21_0_in0(inst_cellmath__19), .inst_cellmath__21_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw2052368036_bdw cynw_cm_float_mul_ieee_I3 (.inst_cellmath__13__1__out0(inst_cellmath__13), .inst_cellmath__13__1__in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw2052368036_bdw cynw_cm_float_mul_ieee_I4 (.inst_cellmath__26__9__out0({N441}), .inst_cellmath__26__9__in0(inst_cellmath__21), .inst_cellmath__26__9__in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I5 (.inst_cellmath__10_0_out0(inst_cellmath__10), .inst_cellmath__10_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw2052368036_bdw cynw_cm_float_mul_ieee_I6 (.inst_cellmath__12__0__out0(inst_cellmath__12), .inst_cellmath__12__0__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I7 (.inst_cellmath__14_0_out0(inst_cellmath__14), .inst_cellmath__14_0_in0(inst_cellmath__12), .inst_cellmath__14_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw2052368036_bdw cynw_cm_float_mul_ieee_I8 (.inst_cellmath__20__3__out0(inst_cellmath__20), .inst_cellmath__20__3__in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw2052368036_bdw cynw_cm_float_mul_ieee_I9 (.inst_cellmath__26__8__out0({N440}), .inst_cellmath__26__8__in0(inst_cellmath__20), .inst_cellmath__26__8__in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I10 (.inst_cellmath__15_0_out0(inst_cellmath__15), .inst_cellmath__15_0_in0(inst_cellmath__12), .inst_cellmath__15_0_in1(inst_cellmath__10));
cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I11 (.inst_cellmath__22_0_out0(inst_cellmath__22), .inst_cellmath__22_0_in0(inst_cellmath__19), .inst_cellmath__22_0_in1(inst_cellmath__17));
cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw2052368036_bdw cynw_cm_float_mul_ieee_I12 (.inst_cellmath__26_1_out0(inst_cellmath__26), .inst_cellmath__26_1_in0({N441}), .inst_cellmath__26_1_in1({N440}), .inst_cellmath__26_1_in2(inst_cellmath__22), .inst_cellmath__26_1_in3(inst_cellmath__15));
cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I13 (.inst_cellmath__23_0_out0(inst_cellmath__23), .inst_cellmath__23_0_in0(b_sign), .inst_cellmath__23_0_in1(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I14 (.inst_cellmath__41_0_out0(x[31]), .inst_cellmath__41_0_in0(inst_cellmath__26), .inst_cellmath__41_0_in1(inst_cellmath__23), .inst_cellmath__41_0_in2(inst_cellmath__22), .inst_cellmath__41_0_in3(inst_cellmath__15), .inst_cellmath__41_0_in4(b_sign), .inst_cellmath__41_0_in5(a_sign));
cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I15 (.inst_cellmath__24_0_out0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}), .inst_cellmath__24_0_in0({b_man[22], b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__24_0_in1({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I16 (.inst_cellmath__25_0_out0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24], inst_cellmath__25[23], inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}), .inst_cellmath__25_0_in0({inst_cellmath__24[47], inst_cellmath__24[46], inst_cellmath__24[45], inst_cellmath__24[44], inst_cellmath__24[43], inst_cellmath__24[42], inst_cellmath__24[41], inst_cellmath__24[40], inst_cellmath__24[39], inst_cellmath__24[38], inst_cellmath__24[37], inst_cellmath__24[36], inst_cellmath__24[35], inst_cellmath__24[34], inst_cellmath__24[33], inst_cellmath__24[32], inst_cellmath__24[31], inst_cellmath__24[30], inst_cellmath__24[29], inst_cellmath__24[28], inst_cellmath__24[27], inst_cellmath__24[26], inst_cellmath__24[25], inst_cellmath__24[24], inst_cellmath__24[23], inst_cellmath__24[22], inst_cellmath__24[21], inst_cellmath__24[20], inst_cellmath__24[19], inst_cellmath__24[18], inst_cellmath__24[17], inst_cellmath__24[16], inst_cellmath__24[15], inst_cellmath__24[14], inst_cellmath__24[13], inst_cellmath__24[12], inst_cellmath__24[11], inst_cellmath__24[10], inst_cellmath__24[9], inst_cellmath__24[8], inst_cellmath__24[7], inst_cellmath__24[6], inst_cellmath__24[5], inst_cellmath__24[4], inst_cellmath__24[3], inst_cellmath__24[2], inst_cellmath__24[1], inst_cellmath__24[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I17 (.inst_cellmath__45_0_out0({inst_cellmath__45[24], inst_cellmath__45[23], inst_cellmath__45[22], inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__45_0_in0({inst_cellmath__25[47], inst_cellmath__25[46], inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw2052368036_bdw cynw_cm_float_mul_ieee_I18 (.inst_cellmath__5_1_out0(inst_cellmath__5), .inst_cellmath__5_1_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw2052368036_bdw cynw_cm_float_mul_ieee_I19 (.inst_cellmath__44__31__out0({N446}), .inst_cellmath__44__31__in0(inst_cellmath__5), .inst_cellmath__44__31__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I20 (.inst_cellmath__6_0_out0(inst_cellmath__6), .inst_cellmath__6_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw2052368036_bdw cynw_cm_float_mul_ieee_I21 (.inst_cellmath__44__30__out0({N445}), .inst_cellmath__44__30__in0(inst_cellmath__6), .inst_cellmath__44__30__in1(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I22 (.inst_cellmath__8_0_out0(inst_cellmath__8), .inst_cellmath__8_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I23 (.inst_cellmath__4_0_out0(inst_cellmath__4), .inst_cellmath__4_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I24 (.inst_cellmath__34_0_out0(inst_cellmath__34), .inst_cellmath__34_0_in0({inst_cellmath__25[22], inst_cellmath__25[21], inst_cellmath__25[20], inst_cellmath__25[19], inst_cellmath__25[18], inst_cellmath__25[17], inst_cellmath__25[16], inst_cellmath__25[15], inst_cellmath__25[14], inst_cellmath__25[13], inst_cellmath__25[12], inst_cellmath__25[11], inst_cellmath__25[10], inst_cellmath__25[9], inst_cellmath__25[8], inst_cellmath__25[7], inst_cellmath__25[6], inst_cellmath__25[5], inst_cellmath__25[4], inst_cellmath__25[3], inst_cellmath__25[2], inst_cellmath__25[1], inst_cellmath__25[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw2052368036_bdw cynw_cm_float_mul_ieee_I25 (.inst_cellmath__44__29__out0({N443}), .inst_cellmath__44__29__in0(inst_cellmath__34), .inst_cellmath__44__29__in1({inst_cellmath__25[24]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw2052368036_bdw cynw_cm_float_mul_ieee_I26 (.inst_cellmath__44__28__out0({N444}), .inst_cellmath__44__28__in0({N443}), .inst_cellmath__44__28__in1(inst_cellmath__4));
cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw2052368036_bdw cynw_cm_float_mul_ieee_I27 (.inst_cellmath__44__27__out0({N447}), .inst_cellmath__44__27__in0(inst_cellmath__8), .inst_cellmath__44__27__in1({N446}), .inst_cellmath__44__27__in2({N445}), .inst_cellmath__44__27__in3({N444}));
cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw2052368036_bdw cynw_cm_float_mul_ieee_I28 (.inst_cellmath__44__26__out0({N448}), .inst_cellmath__44__26__in0({N447}), .inst_cellmath__44__26__in1({inst_cellmath__25[23]}));
cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw2052368036_bdw cynw_cm_float_mul_ieee_I29 (.inst_cellmath__44__33__out0({N449}), .inst_cellmath__44__33__in0({N446}), .inst_cellmath__44__33__in1({N445}));
cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw2052368036_bdw cynw_cm_float_mul_ieee_I30 (.inst_cellmath__44__32__out0({N450}), .inst_cellmath__44__32__in0({N449}), .inst_cellmath__44__32__in1(inst_cellmath__34));
cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I31 (.inst_cellmath__44_0_out0(inst_cellmath__44), .inst_cellmath__44_0_in0({N450}), .inst_cellmath__44_0_in1({N448}));
cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I32 (.inst_cellmath__46_0_out0(inst_cellmath__46), .inst_cellmath__46_0_in0({inst_cellmath__45[24]}), .inst_cellmath__46_0_in1(inst_cellmath__44));
cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I33 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__46), .inst_cellmath__38_0_in1({inst_cellmath__24[47]}));
cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I34 (.inst_cellmath__30_0_out0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}), .inst_cellmath__30_0_in0({b_exp[7], b_exp[6], b_exp[5], b_exp[4], b_exp[3], b_exp[2], b_exp[1], b_exp[0]}), .inst_cellmath__30_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I35 (.inst_cellmath__31_0_out0({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__31_0_in0({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I36 (.inst_cellmath__48_0_out0({inst_cellmath__48[9], inst_cellmath__48[8], inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__48_0_in0(inst_cellmath__38), .inst_cellmath__48_0_in1({inst_cellmath__31[9], inst_cellmath__31[8], inst_cellmath__31[7], inst_cellmath__31[6], inst_cellmath__31[5], inst_cellmath__31[4], inst_cellmath__31[3], inst_cellmath__31[2], inst_cellmath__31[1], inst_cellmath__31[0]}), .inst_cellmath__48_0_in2({inst_cellmath__30[9], inst_cellmath__30[8], inst_cellmath__30[7], inst_cellmath__30[6], inst_cellmath__30[5], inst_cellmath__30[4], inst_cellmath__30[3], inst_cellmath__30[2], inst_cellmath__30[1], inst_cellmath__30[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw2052368036_bdw cynw_cm_float_mul_ieee_I37 (.inst_cellmath__51__49__out0({N461}), .inst_cellmath__51__49__in0({inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw2052368036_bdw cynw_cm_float_mul_ieee_I38 (.inst_cellmath__51__48__out0({N462}), .inst_cellmath__51__48__in0({N461}), .inst_cellmath__51__48__in1({inst_cellmath__48[8]}));
cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I39 (.inst_cellmath__51_0_out0(inst_cellmath__51), .inst_cellmath__51_0_in0({N462}), .inst_cellmath__51_0_in1({inst_cellmath__48[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I40 (.inst_cellmath__28_0_out0(inst_cellmath__28), .inst_cellmath__28_0_in0(inst_cellmath__20), .inst_cellmath__28_0_in1(inst_cellmath__13));
cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I41 (.inst_cellmath__27_0_out0(inst_cellmath__27), .inst_cellmath__27_0_in0(inst_cellmath__21), .inst_cellmath__27_0_in1(inst_cellmath__14));
cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw2052368036_bdw cynw_cm_float_mul_ieee_I42 (.inst_cellmath__50__50__out0({N463}), .inst_cellmath__50__50__in0({inst_cellmath__48[9], inst_cellmath__48[8], inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw2052368036_bdw cynw_cm_float_mul_ieee_I43 (.inst_cellmath__49_1_out0(inst_cellmath__49), .inst_cellmath__49_1_in0(inst_cellmath__51), .inst_cellmath__49_1_in1({N463}), .inst_cellmath__49_1_in2({inst_cellmath__48[9]}), .inst_cellmath__49_1_in3(inst_cellmath__28), .inst_cellmath__49_1_in4(inst_cellmath__27), .inst_cellmath__49_1_in5(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw2052368036_bdw cynw_cm_float_mul_ieee_I44 (.inst_cellmath__37__43__out0({N470}), .inst_cellmath__37__43__in0(inst_cellmath__27), .inst_cellmath__37__43__in1(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw2052368036_bdw cynw_cm_float_mul_ieee_I45 (.inst_cellmath__32__11__out0({N442}), .inst_cellmath__32__11__in0({inst_cellmath__30[8], inst_cellmath__30[7]}));
cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw2052368036_bdw cynw_cm_float_mul_ieee_I46 (.inst_cellmath__32__10__out0(inst_cellmath__32), .inst_cellmath__32__10__in0({N442}), .inst_cellmath__32__10__in1({inst_cellmath__30[9]}));
cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw2052368036_bdw cynw_cm_float_mul_ieee_I47 (.inst_cellmath__37__42__out0({N469}), .inst_cellmath__37__42__in0(inst_cellmath__32), .inst_cellmath__37__42__in1(inst_cellmath__28));
cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I48 (.inst_cellmath__7_0_out0(inst_cellmath__7), .inst_cellmath__7_0_in0({rm[2], rm[1], rm[0]}));
cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I49 (.inst_cellmath__42_0_out0(inst_cellmath__42), .inst_cellmath__42_0_in0(inst_cellmath__7), .inst_cellmath__42_0_in1(inst_cellmath__6), .inst_cellmath__42_0_in2(inst_cellmath__5), .inst_cellmath__42_0_in3(inst_cellmath__23));
cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I50 (.inst_cellmath__52_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__52_0_in0(inst_cellmath__49), .inst_cellmath__52_0_in1({inst_cellmath__48[7], inst_cellmath__48[6], inst_cellmath__48[5], inst_cellmath__48[4], inst_cellmath__48[3], inst_cellmath__48[2], inst_cellmath__48[1], inst_cellmath__48[0]}), .inst_cellmath__52_0_in2(inst_cellmath__42), .inst_cellmath__52_0_in3({N470}), .inst_cellmath__52_0_in4({N469}));
cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw2052368036_bdw cynw_cm_float_mul_ieee_I51 (.inst_cellmath__47_0_out0(inst_cellmath__47), .inst_cellmath__47_0_in0(inst_cellmath__42), .inst_cellmath__47_0_in1(inst_cellmath__32), .inst_cellmath__47_0_in2(inst_cellmath__28), .inst_cellmath__47_0_in3(inst_cellmath__27), .inst_cellmath__47_0_in4(inst_cellmath__26));
cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw2052368036_bdw cynw_cm_float_mul_ieee_I52 (.inst_cellmath__53_U_out0({x[22]}), .inst_cellmath__53_U_in0(inst_cellmath__49), .inst_cellmath__53_U_in1(inst_cellmath__47), .inst_cellmath__53_U_in2({inst_cellmath__45[22]}), .inst_cellmath__53_U_in3(inst_cellmath__44), .inst_cellmath__53_U_in4(inst_cellmath__26), .inst_cellmath__53_U_in5({inst_cellmath__25[46]}));
cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2052368036_bdw cynw_cm_float_mul_ieee_I53 (.inst_cellmath__53_M_out0({x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__53_M_in0(inst_cellmath__49), .inst_cellmath__53_M_in1(inst_cellmath__47), .inst_cellmath__53_M_in2({inst_cellmath__45[21], inst_cellmath__45[20], inst_cellmath__45[19], inst_cellmath__45[18], inst_cellmath__45[17], inst_cellmath__45[16], inst_cellmath__45[15], inst_cellmath__45[14], inst_cellmath__45[13], inst_cellmath__45[12], inst_cellmath__45[11], inst_cellmath__45[10], inst_cellmath__45[9], inst_cellmath__45[8], inst_cellmath__45[7], inst_cellmath__45[6], inst_cellmath__45[5], inst_cellmath__45[4], inst_cellmath__45[3], inst_cellmath__45[2], inst_cellmath__45[1], inst_cellmath__45[0]}), .inst_cellmath__53_M_in3(inst_cellmath__44), .inst_cellmath__53_M_in4(inst_cellmath__26), .inst_cellmath__53_M_in5({inst_cellmath__25[45], inst_cellmath__25[44], inst_cellmath__25[43], inst_cellmath__25[42], inst_cellmath__25[41], inst_cellmath__25[40], inst_cellmath__25[39], inst_cellmath__25[38], inst_cellmath__25[37], inst_cellmath__25[36], inst_cellmath__25[35], inst_cellmath__25[34], inst_cellmath__25[33], inst_cellmath__25[32], inst_cellmath__25[31], inst_cellmath__25[30], inst_cellmath__25[29], inst_cellmath__25[28], inst_cellmath__25[27], inst_cellmath__25[26], inst_cellmath__25[25], inst_cellmath__25[24]}), .inst_cellmath__53_M_in6(inst_cellmath__22), .inst_cellmath__53_M_in7(inst_cellmath__15), .inst_cellmath__53_M_in8({b_man[21], b_man[20], b_man[19], b_man[18], b_man[17], b_man[16], b_man[15], b_man[14], b_man[13], b_man[12], b_man[11], b_man[10], b_man[9], b_man[8], b_man[7], b_man[6], b_man[5], b_man[4], b_man[3], b_man[2], b_man[1], b_man[0]}), .inst_cellmath__53_M_in9({a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__17_0_bdw2052368036_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [7:0] inst_cellmath__17_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__17_0_I0 (.Y(N11), .A(inst_cellmath__17_0_in0[0]), .B(inst_cellmath__17_0_in0[1]));
NAND2XL inst_cellmath__17_0_I1 (.Y(N12), .A(inst_cellmath__17_0_in0[7]), .B(inst_cellmath__17_0_in0[6]));
NAND2XL inst_cellmath__17_0_I2 (.Y(N13), .A(inst_cellmath__17_0_in0[5]), .B(inst_cellmath__17_0_in0[4]));
NAND2XL inst_cellmath__17_0_I3 (.Y(N14), .A(inst_cellmath__17_0_in0[3]), .B(inst_cellmath__17_0_in0[2]));
NOR2XL inst_cellmath__17_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__17_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__17_0_I6 (.Y(inst_cellmath__17_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__19__2__bdw2052368036_bdw (
	inst_cellmath__19__2__out0,
	inst_cellmath__19__2__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__19__2__out0;
input [22:0] inst_cellmath__19__2__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__19__2__I1 (.Y(N27), .A(inst_cellmath__19__2__in0[22]), .B(inst_cellmath__19__2__in0[21]));
NOR2XL inst_cellmath__19__2__I2 (.Y(N28), .A(inst_cellmath__19__2__in0[20]), .B(inst_cellmath__19__2__in0[19]));
NOR2XL inst_cellmath__19__2__I3 (.Y(N29), .A(inst_cellmath__19__2__in0[18]), .B(inst_cellmath__19__2__in0[17]));
NOR2XL inst_cellmath__19__2__I4 (.Y(N30), .A(inst_cellmath__19__2__in0[16]), .B(inst_cellmath__19__2__in0[15]));
NOR2XL inst_cellmath__19__2__I5 (.Y(N31), .A(inst_cellmath__19__2__in0[14]), .B(inst_cellmath__19__2__in0[13]));
NOR2XL inst_cellmath__19__2__I6 (.Y(N32), .A(inst_cellmath__19__2__in0[12]), .B(inst_cellmath__19__2__in0[11]));
NOR2XL inst_cellmath__19__2__I7 (.Y(N33), .A(inst_cellmath__19__2__in0[10]), .B(inst_cellmath__19__2__in0[9]));
NOR2XL inst_cellmath__19__2__I8 (.Y(N34), .A(inst_cellmath__19__2__in0[8]), .B(inst_cellmath__19__2__in0[7]));
NOR2XL inst_cellmath__19__2__I9 (.Y(N35), .A(inst_cellmath__19__2__in0[6]), .B(inst_cellmath__19__2__in0[5]));
NOR2XL inst_cellmath__19__2__I10 (.Y(N36), .A(inst_cellmath__19__2__in0[4]), .B(inst_cellmath__19__2__in0[3]));
NAND2XL inst_cellmath__19__2__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__19__2__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__19__2__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__19__2__I25 (.Y(N44), .A(inst_cellmath__19__2__in0[0]), .B(inst_cellmath__19__2__in0[1]), .C(inst_cellmath__19__2__in0[2]), .D(N39));
NOR2XL inst_cellmath__19__2__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__19__2__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__19__2__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__19__2__I23 (.Y(inst_cellmath__19__2__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__21_0_bdw2052368036_bdw (
	inst_cellmath__21_0_out0,
	inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__21_0_out0;
input  inst_cellmath__21_0_in0,
	inst_cellmath__21_0_in1;
AND2XL inst_cellmath__21_0_I0 (.Y(inst_cellmath__21_0_out0), .A(inst_cellmath__21_0_in1), .B(inst_cellmath__21_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__13__1__bdw2052368036_bdw (
	inst_cellmath__13__1__out0,
	inst_cellmath__13__1__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__13__1__out0;
input [7:0] inst_cellmath__13__1__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__13__1__I0 (.Y(N11), .A(inst_cellmath__13__1__in0[0]), .B(inst_cellmath__13__1__in0[1]));
NOR2XL inst_cellmath__13__1__I1 (.Y(N12), .A(inst_cellmath__13__1__in0[7]), .B(inst_cellmath__13__1__in0[6]));
NOR2XL inst_cellmath__13__1__I2 (.Y(N13), .A(inst_cellmath__13__1__in0[5]), .B(inst_cellmath__13__1__in0[4]));
NOR2XL inst_cellmath__13__1__I3 (.Y(N14), .A(inst_cellmath__13__1__in0[3]), .B(inst_cellmath__13__1__in0[2]));
NAND2XL inst_cellmath__13__1__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__13__1__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__13__1__I6 (.Y(inst_cellmath__13__1__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__9__bdw2052368036_bdw (
	inst_cellmath__26__9__out0,
	inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__9__out0;
input  inst_cellmath__26__9__in0,
	inst_cellmath__26__9__in1;
AND2XL inst_cellmath__26__9__I0 (.Y(inst_cellmath__26__9__out0[0]), .A(inst_cellmath__26__9__in1), .B(inst_cellmath__26__9__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__10_0_bdw2052368036_bdw (
	inst_cellmath__10_0_out0,
	inst_cellmath__10_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__10_0_out0;
input [7:0] inst_cellmath__10_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__10_0_I0 (.Y(N11), .A(inst_cellmath__10_0_in0[0]), .B(inst_cellmath__10_0_in0[1]));
NAND2XL inst_cellmath__10_0_I1 (.Y(N12), .A(inst_cellmath__10_0_in0[7]), .B(inst_cellmath__10_0_in0[6]));
NAND2XL inst_cellmath__10_0_I2 (.Y(N13), .A(inst_cellmath__10_0_in0[5]), .B(inst_cellmath__10_0_in0[4]));
NAND2XL inst_cellmath__10_0_I3 (.Y(N14), .A(inst_cellmath__10_0_in0[3]), .B(inst_cellmath__10_0_in0[2]));
NOR2XL inst_cellmath__10_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__10_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__10_0_I6 (.Y(inst_cellmath__10_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__12__0__bdw2052368036_bdw (
	inst_cellmath__12__0__out0,
	inst_cellmath__12__0__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__12__0__out0;
input [22:0] inst_cellmath__12__0__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__12__0__I1 (.Y(N27), .A(inst_cellmath__12__0__in0[22]), .B(inst_cellmath__12__0__in0[21]));
NOR2XL inst_cellmath__12__0__I2 (.Y(N28), .A(inst_cellmath__12__0__in0[20]), .B(inst_cellmath__12__0__in0[19]));
NOR2XL inst_cellmath__12__0__I3 (.Y(N29), .A(inst_cellmath__12__0__in0[18]), .B(inst_cellmath__12__0__in0[17]));
NOR2XL inst_cellmath__12__0__I4 (.Y(N30), .A(inst_cellmath__12__0__in0[16]), .B(inst_cellmath__12__0__in0[15]));
NOR2XL inst_cellmath__12__0__I5 (.Y(N31), .A(inst_cellmath__12__0__in0[14]), .B(inst_cellmath__12__0__in0[13]));
NOR2XL inst_cellmath__12__0__I6 (.Y(N32), .A(inst_cellmath__12__0__in0[12]), .B(inst_cellmath__12__0__in0[11]));
NOR2XL inst_cellmath__12__0__I7 (.Y(N33), .A(inst_cellmath__12__0__in0[10]), .B(inst_cellmath__12__0__in0[9]));
NOR2XL inst_cellmath__12__0__I8 (.Y(N34), .A(inst_cellmath__12__0__in0[8]), .B(inst_cellmath__12__0__in0[7]));
NOR2XL inst_cellmath__12__0__I9 (.Y(N35), .A(inst_cellmath__12__0__in0[6]), .B(inst_cellmath__12__0__in0[5]));
NOR2XL inst_cellmath__12__0__I10 (.Y(N36), .A(inst_cellmath__12__0__in0[4]), .B(inst_cellmath__12__0__in0[3]));
NAND2XL inst_cellmath__12__0__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__12__0__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__12__0__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__12__0__I25 (.Y(N44), .A(inst_cellmath__12__0__in0[0]), .B(inst_cellmath__12__0__in0[1]), .C(inst_cellmath__12__0__in0[2]), .D(N39));
NOR2XL inst_cellmath__12__0__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__12__0__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__12__0__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__12__0__I23 (.Y(inst_cellmath__12__0__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__14_0_bdw2052368036_bdw (
	inst_cellmath__14_0_out0,
	inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__14_0_out0;
input  inst_cellmath__14_0_in0,
	inst_cellmath__14_0_in1;
AND2XL inst_cellmath__14_0_I0 (.Y(inst_cellmath__14_0_out0), .A(inst_cellmath__14_0_in1), .B(inst_cellmath__14_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__20__3__bdw2052368036_bdw (
	inst_cellmath__20__3__out0,
	inst_cellmath__20__3__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__20__3__out0;
input [7:0] inst_cellmath__20__3__in0;
wire N11,N12,N13,N14,N15,N16;
NOR2XL inst_cellmath__20__3__I0 (.Y(N11), .A(inst_cellmath__20__3__in0[0]), .B(inst_cellmath__20__3__in0[1]));
NOR2XL inst_cellmath__20__3__I1 (.Y(N12), .A(inst_cellmath__20__3__in0[7]), .B(inst_cellmath__20__3__in0[6]));
NOR2XL inst_cellmath__20__3__I2 (.Y(N13), .A(inst_cellmath__20__3__in0[5]), .B(inst_cellmath__20__3__in0[4]));
NOR2XL inst_cellmath__20__3__I3 (.Y(N14), .A(inst_cellmath__20__3__in0[3]), .B(inst_cellmath__20__3__in0[2]));
NAND2XL inst_cellmath__20__3__I4 (.Y(N15), .A(N11), .B(N12));
NAND2XL inst_cellmath__20__3__I5 (.Y(N16), .A(N13), .B(N14));
NOR2XL inst_cellmath__20__3__I6 (.Y(inst_cellmath__20__3__out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26__8__bdw2052368036_bdw (
	inst_cellmath__26__8__out0,
	inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__26__8__out0;
input  inst_cellmath__26__8__in0,
	inst_cellmath__26__8__in1;
AND2XL inst_cellmath__26__8__I0 (.Y(inst_cellmath__26__8__out0[0]), .A(inst_cellmath__26__8__in0), .B(inst_cellmath__26__8__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__15_0_bdw2052368036_bdw (
	inst_cellmath__15_0_out0,
	inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__15_0_out0;
input  inst_cellmath__15_0_in0,
	inst_cellmath__15_0_in1;
NOR2BX1 inst_cellmath__15_0_I2 (.Y(inst_cellmath__15_0_out0), .AN(inst_cellmath__15_0_in1), .B(inst_cellmath__15_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__22_0_bdw2052368036_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__22_0_out0;
input  inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1;
NOR2BX1 inst_cellmath__22_0_I2 (.Y(inst_cellmath__22_0_out0), .AN(inst_cellmath__22_0_in1), .B(inst_cellmath__22_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__26_1_bdw2052368036_bdw (
	inst_cellmath__26_1_out0,
	inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1,
	inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__26_1_out0;
input [0:0] inst_cellmath__26_1_in0,
	inst_cellmath__26_1_in1;
input  inst_cellmath__26_1_in2,
	inst_cellmath__26_1_in3;
OR4X1 inst_cellmath__26_1_I6 (.Y(inst_cellmath__26_1_out0), .A(inst_cellmath__26_1_in2), .B(inst_cellmath__26_1_in3), .C(inst_cellmath__26_1_in0[0]), .D(inst_cellmath__26_1_in1[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__23_0_bdw2052368036_bdw (
	inst_cellmath__23_0_out0,
	inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__23_0_out0;
input  inst_cellmath__23_0_in0,
	inst_cellmath__23_0_in1;
XOR2XL inst_cellmath__23_0_I0 (.Y(inst_cellmath__23_0_out0), .A(inst_cellmath__23_0_in1), .B(inst_cellmath__23_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__41_0_bdw2052368036_bdw (
	inst_cellmath__41_0_out0,
	inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__41_0_out0;
input  inst_cellmath__41_0_in0,
	inst_cellmath__41_0_in1,
	inst_cellmath__41_0_in2,
	inst_cellmath__41_0_in3,
	inst_cellmath__41_0_in4,
	inst_cellmath__41_0_in5;
wire N14,N16;
NAND2BXL inst_cellmath__41_0_I6 (.Y(N14), .AN(inst_cellmath__41_0_in4), .B(inst_cellmath__41_0_in2));
MX2XL inst_cellmath__41_0_I3 (.Y(N16), .A(N14), .B(inst_cellmath__41_0_in5), .S0(inst_cellmath__41_0_in3));
MX2XL inst_cellmath__41_0_I5 (.Y(inst_cellmath__41_0_out0), .A(inst_cellmath__41_0_in1), .B(N16), .S0(inst_cellmath__41_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__24_0_bdw2052368036_bdw (
	inst_cellmath__24_0_out0,
	inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__24_0_out0;
input [22:0] inst_cellmath__24_0_in0,
	inst_cellmath__24_0_in1;
wire N372,N373,N381,N382,N384,N385,N386 
	,N387,N388,N389,N390,N391,N392,N393,N394 
	,N395,N396,N397,N398,N399,N400,N401,N402 
	,N403,N404,N405,N406,N407,N408,N409,N410 
	,N411,N412,N413,N414,N415,N416,N417,N418 
	,N419,N420,N421,N422,N423,N424,N425,N426 
	,N427,N428,N429,N433,N438,N439,N443,N444 
	,N445,N446,N447,N448,N449,N450,N451,N452 
	,N453,N454,N455,N456,N457,N458,N459,N460 
	,N461,N462,N463,N464,N465,N466,N467,N468 
	,N469,N470,N471,N472,N473,N474,N475,N476 
	,N477,N478,N479,N480,N481,N482,N483,N484 
	,N485,N486,N487,N488,N489,N490,N491,N492 
	,N493,N497,N502,N503,N507,N508,N509,N510 
	,N511,N512,N513,N514,N515,N516,N517,N518 
	,N519,N520,N521,N522,N523,N524,N525,N526 
	,N527,N528,N529,N530,N531,N532,N533,N534 
	,N535,N536,N537,N538,N539,N540,N541,N542 
	,N543,N544,N545,N546,N547,N548,N549,N550 
	,N551,N552,N553,N554,N555,N556,N557,N561 
	,N566,N567,N571,N572,N573,N574,N575,N576 
	,N577,N578,N579,N580,N581,N582,N583,N584 
	,N585,N586,N587,N588,N589,N590,N591,N592 
	,N593,N594,N595,N596,N597,N598,N599,N600 
	,N601,N602,N603,N604,N605,N606,N607,N608 
	,N609,N610,N611,N612,N613,N614,N615,N616 
	,N617,N618,N619,N620,N621,N625,N630,N631 
	,N635,N636,N637,N638,N639,N640,N641,N642 
	,N643,N644,N645,N646,N647,N648,N649,N650 
	,N651,N652,N653,N654,N655,N656,N657,N658 
	,N659,N660,N661,N662,N663,N664,N665,N666 
	,N667,N668,N669,N670,N671,N672,N673,N674 
	,N675,N676,N677,N678,N679,N680,N681,N682 
	,N683,N684,N685,N689,N694,N695,N699,N700 
	,N701,N702,N703,N704,N705,N706,N707,N708 
	,N709,N710,N711,N712,N713,N714,N715,N716 
	,N717,N718,N719,N720,N721,N722,N723,N724 
	,N725,N726,N727,N728,N729,N730,N731,N732 
	,N733,N734,N735,N736,N737,N738,N739,N740 
	,N741,N742,N743,N744,N745,N746,N747,N748 
	,N749,N753,N758,N759,N763,N764,N765,N766 
	,N767,N768,N769,N770,N771,N772,N773,N774 
	,N775,N776,N777,N778,N779,N780,N781,N782 
	,N783,N784,N785,N786,N787,N788,N789,N790 
	,N791,N792,N793,N794,N795,N796,N797,N798 
	,N799,N800,N801,N802,N803,N804,N805,N806 
	,N807,N808,N809,N810,N811,N812,N813,N817 
	,N822,N823,N827,N828,N829,N830,N831,N832 
	,N833,N834,N835,N836,N837,N838,N839,N840 
	,N841,N842,N843,N844,N845,N846,N847,N848 
	,N849,N850,N851,N852,N853,N854,N855,N856 
	,N857,N858,N859,N860,N861,N862,N863,N864 
	,N865,N866,N867,N868,N869,N870,N871,N872 
	,N873,N874,N875,N876,N877,N881,N886,N887 
	,N891,N892,N893,N894,N895,N896,N897,N898 
	,N899,N900,N901,N902,N903,N904,N905,N906 
	,N907,N908,N909,N910,N911,N912,N913,N914 
	,N915,N916,N917,N918,N919,N920,N921,N922 
	,N923,N924,N925,N926,N927,N928,N929,N930 
	,N931,N932,N933,N934,N935,N936,N937,N938 
	,N939,N940,N941,N945,N950,N951,N955,N956 
	,N957,N958,N959,N960,N961,N962,N963,N964 
	,N965,N966,N967,N968,N969,N970,N971,N972 
	,N973,N974,N975,N976,N977,N978,N979,N980 
	,N981,N982,N983,N984,N985,N986,N987,N988 
	,N989,N990,N991,N992,N993,N994,N995,N996 
	,N997,N998,N999,N1000,N1001,N1002,N1003,N1004 
	,N1005,N1009,N1014,N1015,N1019,N1020,N1021,N1022 
	,N1023,N1024,N1025,N1026,N1027,N1028,N1029,N1030 
	,N1031,N1032,N1033,N1034,N1035,N1036,N1037,N1038 
	,N1039,N1040,N1041,N1042,N1043,N1044,N1045,N1046 
	,N1047,N1048,N1049,N1050,N1051,N1052,N1053,N1054 
	,N1055,N1056,N1057,N1058,N1059,N1060,N1061,N1062 
	,N1063,N1064,N1065,N1066,N1067,N1068,N1069,N1073 
	,N1078,N1084,N1092,N1093,N1094,N1095,N1096,N1097 
	,N1098,N1099,N1100,N1101,N1102,N1103,N1104,N1105 
	,N1106,N1107,N1108,N1109,N1110,N1111,N1112,N1113 
	,N1114,N1115,N1116,N1117,N1118,N1119,N1120,N1121 
	,N1122,N1123,N1124,N1125,N1126,N1127,N1128,N1129 
	,N1130,N1131,N1132,N1133,N1134,N1135,N1136,N1137 
	,N1138,N1140,N1144,N1212,N1213,N1214,N1215,N1216 
	,N1217,N1218,N1219,N1220,N1221,N1222,N1223,N1224 
	,N1225,N1226,N1227,N1228,N1229,N1230,N1231,N1232 
	,N1233,N1234,N1235,N1236,N1237,N1238,N1239,N1240 
	,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248 
	,N1249,N1250,N1251,N1252,N1253,N1254,N1255,N1256 
	,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264 
	,N1265,N1266,N1267,N1268,N1269,N1270,N1271,N1272 
	,N1273,N1274,N1275,N1276,N1277,N1278,N1279,N1280 
	,N1281,N1282,N1283,N1284,N1285,N1286,N1287,N1288 
	,N1289,N1290,N1291,N1292,N1293,N1294,N1295,N1296 
	,N1297,N1298,N1299,N1300,N1301,N1302,N1303,N1304 
	,N1305,N1306,N1307,N1308,N1309,N1310,N1311,N1312 
	,N1313,N1314,N1315,N1316,N1317,N1318,N1319,N1320 
	,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328 
	,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336 
	,N1337,N1338,N1339,N1340,N1341,N1342,N1343,N1344 
	,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352 
	,N1353,N1354,N1355,N1356,N1357,N1358,N1359,N1360 
	,N1361,N1362,N1363,N1364,N1365,N1366,N1367,N1368 
	,N1369,N1370,N1371,N1372,N1373,N1374,N1375,N1376 
	,N1377,N1378,N1379,N1380,N1381,N1382,N1383,N1384 
	,N1385,N1386,N1387,N1388,N1389,N1390,N1391,N1392 
	,N1393,N1394,N1395,N1396,N1397,N1398,N1399,N1400 
	,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408 
	,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416 
	,N1417,N1418,N1419,N1420,N1421,N1422,N1423,N1424 
	,N1425,N1426,N1427,N1428,N1429,N1430,N1431,N1432 
	,N1433,N1434,N1435,N1436,N1437,N1438,N1439,N1440 
	,N1441,N1442,N1443,N1444,N1445,N1446,N1447,N1448 
	,N1449,N1450,N1451,N1452,N1453,N1454,N1455,N1458 
	,N1459,N1460,N1461,N1462,N1463,N1464,N1465,N1466 
	,N1467,N1468,N1469,N1470,N1471,N1472,N1473,N1474 
	,N1477,N1478,N1479,N1480,N1481,N1482,N1483,N1484 
	,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492 
	,N1493,N1494,N1495,N1496,N1497,N1498,N1499,N1500 
	,N1501,N1502,N1503,N1504,N1505,N1506,N1507,N1508 
	,N1509,N1510,N1513,N1514,N1515,N1516,N1517,N1518 
	,N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526 
	,N1527,N1528,N1529,N1530,N1531,N1532,N1533,N1534 
	,N1535,N1536,N1537,N1538,N1539,N1540,N1541,N1542 
	,N1543,N1546,N1547,N1548,N1549,N1550,N1551,N1552 
	,N1553,N1554,N1555,N1556,N1557,N1558,N1559,N1560 
	,N1561,N1562,N1563,N1564,N1565,N1566,N1567,N1568 
	,N1569,N1570,N1571,N1572,N1573,N1576,N1577,N1578 
	,N1579,N1580,N1581,N1582,N1583,N1584,N1585,N1586 
	,N1587,N1588,N1589,N1590,N1591,N1592,N1593,N1594 
	,N1595,N1596,N1597,N1598,N1599,N1600,N1603,N1604 
	,N1605,N1606,N1607,N1608,N1609,N1610,N1611,N1612 
	,N1613,N1614,N1615,N1616,N1617,N1618,N1619,N1620 
	,N1621,N1622,N1623,N1624,N1627,N1628,N1629,N1630 
	,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638 
	,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1648 
	,N1649,N1650,N1651,N1652,N1653,N1654,N1655,N1656 
	,N1657,N1658,N1659,N1660,N1661,N1662,N1663,N1666 
	,N1667,N1668,N1669,N1670,N1671,N1672,N1673,N1674 
	,N1675,N1676,N1677,N1678,N1681,N1682,N1683,N1684 
	,N1685,N1686,N1687,N1688,N1689,N1690,N1693,N1694 
	,N1695,N1696,N1697,N1702,N1703,N1708,N1710,N1712 
	,N1713,N1714,N1715,N1716,N1717,N1718,N1719,N1720 
	,N1721,N1722,N1723,N1724,N1725,N1726,N1727,N1728 
	,N1729,N1730,N1731,N1732,N1733,N1734,N1735,N1736 
	,N1737,N1738,N1739,N1740,N1741,N1742,N1743,N1744 
	,N1745,N1748,N1758,N1766,N1778,N1790,N1806,N1822 
	,N1842,N1862,N1866,N1867,N1890,N1924,N1926,N1930 
	,N1931,N1962,N1966,N1967,N1974,N1975,N2008,N2010 
	,N2042,N2045,N2048,N2051,N2054,N2057,N2060,N2063 
	,N2066,N2069,N2072,N2075,N2078,N2081,N2084,N2087 
	,N2090,N2110,N2113,N2114,N2115,N2116,N2117,N2118 
	,N2119,N2120,N2121,N2122,N2123,N2124,N2125,N2126 
	,N2127,N2128,N2129,N2130,N2131,N2132,N2133,N2134 
	,N2135,N2136,N2137,N2138,N2139,N2140,N2141,N2142 
	,N2143,N2144,N2145,N2146,N2147,N2148,N2149,N2150 
	,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158 
	,N2159,N2160,N2161,N2162,N2163,N2164,N2165,N2166 
	,N2167,N2169,N2170,N2172,N2173,N2174,N2175,N2176 
	,N2177,N2178,N2179,N2180,N2181,N2182,N2183,N2184 
	,N2185,N2186,N2187,N2188,N2189,N2190,N2191,N2192 
	,N2193,N2194,N2195,N2196,N2197,N2200,N2202,N2203 
	,N2204,N2205,N2206,N2207,N2208,N2209,N2210,N2211 
	,N2214,N2216,N2217,N2218,N2220,N2222,N2223,N2224 
	,N2228,N2231,N2232,N2234,N2235,N2236,N2240,N2244 
	,N2245,N2246,N2250,N2254,N2258,N2261,N2262,N2264 
	,N2265,N2266,N2270,N2274,N2275,N2276,N2280,N2284 
	,N2288,N2289,N2290,N2294,N2295,N2296,N2300,N2304 
	,N2308,N2312,N2316,N2320,N2324,N2737,N2964,N3191 
	,N3418,N3645,N3872,N4099,N4326,N4553,N4780,N5216 
	,N5229,N5242,N5255,N5268,N5281,N5294,N5307,N5320 
	,N5333,N5346,N5359,N5372,N5385,N5398,N5411,N5424 
	,N5437,N5450,N5463,N5476,N5489,N5502,N5515,N5528 
	,N5541,N5554,N5567,N5580,N5593,N5606,N5619,N5632 
	,N5645,N5658,N5671,N5684,N5697,N5710,N5723,N5736 
	,N5749,N5762,N5775,N5788,N5801,N5814,N5827,N5840 
	,N5853,N5866,N5879,N5892,N5905,N5918,N5935,N5940 
	,N5953,N5966,N5979,N5992,N6009,N6014,N6027,N6040 
	,N6053,N6066,N6079,N6092,N6105,N6118,N6131,N6148 
	,N6153,N6166,N6179,N6192,N6205,N6218,N6231,N6244 
	,N6257,N6274,N6279,N6292,N6305,N6318,N6331,N6344 
	,N6357,N6370,N6387,N6392,N6405,N6418,N6431,N6444 
	,N6457,N6470,N6487,N6492,N6505,N6518,N6531,N6544 
	,N6557,N6574,N6579,N6592,N6605,N6618,N6631,N6648 
	,N6653,N6666,N6679,N6692,N6709,N6714,N6727,N6740 
	,N6757,N6762,N6775,N6792,N6797,N6909,N6910,N6911 
	,N6912,N6913,N6914,N6915,N6916,N6917,N6918,N6919 
	,N6920,N6921,N6922,N6923,N6924,N6925,N6926,N6927 
	,N6928,N6929,N6930,N6931,N6936,N6937,N6942,N6947 
	,N6952,N6957,N6962,N6967,N6972,N6977,N6982,N6987 
	,N6990,N6991,N6992,N6999,N7000,N7010,N7011,N7025 
	,N7026,N7064,N7100,N7101,N7104,N7105,N7116,N7120 
	,N7128,N7131,N7132,N7133,N7134,N7135,N7162,N7169 
	;
INVXL inst_cellmath__24_0_I2258 (.Y(N6909), .A(inst_cellmath__24_0_in1[0]));
INVXL inst_cellmath__24_0_I2259 (.Y(N6910), .A(inst_cellmath__24_0_in1[1]));
INVXL inst_cellmath__24_0_I2260 (.Y(N6911), .A(inst_cellmath__24_0_in1[2]));
INVXL inst_cellmath__24_0_I2261 (.Y(N6912), .A(inst_cellmath__24_0_in1[3]));
INVXL inst_cellmath__24_0_I2262 (.Y(N6913), .A(inst_cellmath__24_0_in1[4]));
INVXL inst_cellmath__24_0_I2263 (.Y(N6914), .A(inst_cellmath__24_0_in1[5]));
INVXL inst_cellmath__24_0_I2264 (.Y(N6915), .A(inst_cellmath__24_0_in1[6]));
INVXL inst_cellmath__24_0_I2265 (.Y(N6916), .A(inst_cellmath__24_0_in1[7]));
INVXL inst_cellmath__24_0_I2266 (.Y(N6917), .A(inst_cellmath__24_0_in1[8]));
INVXL inst_cellmath__24_0_I2267 (.Y(N6918), .A(inst_cellmath__24_0_in1[9]));
INVXL inst_cellmath__24_0_I2268 (.Y(N6919), .A(inst_cellmath__24_0_in1[10]));
INVXL inst_cellmath__24_0_I2269 (.Y(N6920), .A(inst_cellmath__24_0_in1[11]));
INVXL inst_cellmath__24_0_I2270 (.Y(N6921), .A(inst_cellmath__24_0_in1[12]));
INVXL inst_cellmath__24_0_I2271 (.Y(N6922), .A(inst_cellmath__24_0_in1[13]));
INVXL inst_cellmath__24_0_I2272 (.Y(N6923), .A(inst_cellmath__24_0_in1[14]));
INVXL inst_cellmath__24_0_I2273 (.Y(N6924), .A(inst_cellmath__24_0_in1[15]));
INVXL inst_cellmath__24_0_I2274 (.Y(N6925), .A(inst_cellmath__24_0_in1[16]));
INVXL inst_cellmath__24_0_I2275 (.Y(N6926), .A(inst_cellmath__24_0_in1[17]));
INVXL inst_cellmath__24_0_I2276 (.Y(N6927), .A(inst_cellmath__24_0_in1[18]));
INVXL inst_cellmath__24_0_I2277 (.Y(N6928), .A(inst_cellmath__24_0_in1[19]));
INVXL inst_cellmath__24_0_I2278 (.Y(N6929), .A(inst_cellmath__24_0_in1[20]));
INVXL inst_cellmath__24_0_I2279 (.Y(N6930), .A(inst_cellmath__24_0_in1[21]));
INVXL inst_cellmath__24_0_I2280 (.Y(N6931), .A(inst_cellmath__24_0_in1[22]));
INVXL enc3_A_I1368 (.Y(N372), .A(inst_cellmath__24_0_in0[0]));
NAND2X1 enc3_A_I1371 (.Y(N373), .A(inst_cellmath__24_0_in0[1]), .B(N372));
INVXL inst_cellmath__24_0_I2285 (.Y(N6936), .A(inst_cellmath__24_0_in0[1]));
XNOR2X1 addgen4_A_I1372 (.Y(N382), .A(N6909), .B(N6936));
OAI22XL addgen4_A_I1373 (.Y(N381), .A0(N382), .A1(N372), .B0(N6936), .B1(N373));
XNOR2X1 inst_cellmath__24_0_I1374 (.Y(N384), .A(N6910), .B(N6936));
OA22X1 inst_cellmath__24_0_I2510 (.Y(N6937), .A0(N384), .A1(N372), .B0(N382), .B1(N373));
XNOR2X1 addgen4_A_I1376 (.Y(N386), .A(N6911), .B(N6936));
OAI22XL addgen4_A_I1377 (.Y(N385), .A0(N386), .A1(N372), .B0(N384), .B1(N373));
XNOR2X1 addgen4_A_I1378 (.Y(N388), .A(N6912), .B(N6936));
OAI22XL addgen4_A_I1379 (.Y(N387), .A0(N388), .A1(N372), .B0(N386), .B1(N373));
XNOR2X1 addgen4_A_I1380 (.Y(N390), .A(N6913), .B(N6936));
OAI22XL addgen4_A_I1381 (.Y(N389), .A0(N390), .A1(N372), .B0(N388), .B1(N373));
XNOR2X1 addgen4_A_I1382 (.Y(N392), .A(N6914), .B(N6936));
OAI22XL addgen4_A_I1383 (.Y(N391), .A0(N392), .A1(N372), .B0(N390), .B1(N373));
XNOR2X1 addgen4_A_I1384 (.Y(N394), .A(N6915), .B(N6936));
OAI22XL addgen4_A_I1385 (.Y(N393), .A0(N394), .A1(N372), .B0(N392), .B1(N373));
XNOR2X1 addgen4_A_I1386 (.Y(N396), .A(N6916), .B(N6936));
OAI22XL addgen4_A_I1387 (.Y(N395), .A0(N396), .A1(N372), .B0(N394), .B1(N373));
XNOR2X1 addgen4_A_I1388 (.Y(N398), .A(N6917), .B(N6936));
OAI22XL addgen4_A_I1389 (.Y(N397), .A0(N398), .A1(N372), .B0(N396), .B1(N373));
XNOR2X1 addgen4_A_I1390 (.Y(N400), .A(N6918), .B(N6936));
OAI22XL addgen4_A_I1391 (.Y(N399), .A0(N400), .A1(N372), .B0(N398), .B1(N373));
XNOR2X1 addgen4_A_I1392 (.Y(N402), .A(N6919), .B(N6936));
OAI22XL addgen4_A_I1393 (.Y(N401), .A0(N402), .A1(N372), .B0(N400), .B1(N373));
XNOR2X1 addgen4_A_I1394 (.Y(N404), .A(N6920), .B(N6936));
OAI22XL addgen4_A_I1395 (.Y(N403), .A0(N404), .A1(N372), .B0(N402), .B1(N373));
XNOR2X1 addgen4_A_I1396 (.Y(N406), .A(N6921), .B(N6936));
OAI22XL addgen4_A_I1397 (.Y(N405), .A0(N406), .A1(N372), .B0(N404), .B1(N373));
XNOR2X1 addgen4_A_I1398 (.Y(N408), .A(N6922), .B(N6936));
OAI22XL addgen4_A_I1399 (.Y(N407), .A0(N408), .A1(N372), .B0(N406), .B1(N373));
XNOR2X1 addgen4_A_I1400 (.Y(N410), .A(N6923), .B(N6936));
OAI22XL addgen4_A_I1401 (.Y(N409), .A0(N410), .A1(N372), .B0(N408), .B1(N373));
XNOR2X1 addgen4_A_I1402 (.Y(N412), .A(N6924), .B(N6936));
OAI22XL addgen4_A_I1403 (.Y(N411), .A0(N412), .A1(N372), .B0(N410), .B1(N373));
XNOR2X1 addgen4_A_I1404 (.Y(N414), .A(N6925), .B(N6936));
OAI22XL addgen4_A_I1405 (.Y(N413), .A0(N414), .A1(N372), .B0(N412), .B1(N373));
XNOR2X1 addgen4_A_I1406 (.Y(N416), .A(N6926), .B(N6936));
OAI22XL addgen4_A_I1407 (.Y(N415), .A0(N416), .A1(N372), .B0(N414), .B1(N373));
XNOR2X1 addgen4_A_I1408 (.Y(N418), .A(N6927), .B(N6936));
OAI22XL addgen4_A_I1409 (.Y(N417), .A0(N418), .A1(N372), .B0(N416), .B1(N373));
XNOR2X1 addgen4_A_I1410 (.Y(N420), .A(N6928), .B(N6936));
OAI22XL addgen4_A_I1411 (.Y(N419), .A0(N420), .A1(N372), .B0(N418), .B1(N373));
XNOR2X1 addgen4_A_I1412 (.Y(N422), .A(N6929), .B(N6936));
OAI22XL addgen4_A_I1413 (.Y(N421), .A0(N422), .A1(N372), .B0(N420), .B1(N373));
XNOR2X1 addgen4_A_I1414 (.Y(N424), .A(N6930), .B(N6936));
OAI22XL addgen4_A_I1415 (.Y(N423), .A0(N424), .A1(N372), .B0(N422), .B1(N373));
XNOR2X1 addgen4_A_I1416 (.Y(N426), .A(N6931), .B(N6936));
OAI22XL addgen4_A_I1417 (.Y(N425), .A0(N426), .A1(N372), .B0(N424), .B1(N373));
INVXL addgen4_A_I1418 (.Y(N428), .A(N6936));
OAI22XL addgen4_A_I1419 (.Y(N427), .A0(N428), .A1(N372), .B0(N426), .B1(N373));
MXI2XL inst_cellmath__24_0_I113 (.Y(N429), .A(N373), .B(N372), .S0(N428));
AOI21XL inst_cellmath__24_0_I114 (.Y(N433), .A0(N372), .A1(N373), .B0(N6936));
XNOR2X1 enc3_A_I1420 (.Y(N438), .A(inst_cellmath__24_0_in0[2]), .B(inst_cellmath__24_0_in0[1]));
XOR2XL enc3_A_I1421 (.Y(N2737), .A(inst_cellmath__24_0_in0[3]), .B(inst_cellmath__24_0_in0[1]));
NAND2X1 enc3_A_I1423 (.Y(N439), .A(N2737), .B(N438));
INVXL inst_cellmath__24_0_I2291 (.Y(N6942), .A(inst_cellmath__24_0_in0[3]));
NAND2XL inst_cellmath__24_0_I119 (.Y(N443), .A(inst_cellmath__24_0_in0[1]), .B(inst_cellmath__24_0_in0[2]));
AND2XL inst_cellmath__24_0_I120 (.Y(N444), .A(inst_cellmath__24_0_in0[3]), .B(N443));
XNOR2X1 addgen4_A_I1424 (.Y(N446), .A(N6909), .B(N6942));
OAI22XL addgen4_A_I1425 (.Y(N445), .A0(N446), .A1(N438), .B0(N6942), .B1(N439));
XNOR2X1 addgen4_A_I1426 (.Y(N448), .A(N6910), .B(N6942));
OAI22XL addgen4_A_I1427 (.Y(N447), .A0(N448), .A1(N438), .B0(N446), .B1(N439));
XNOR2X1 addgen4_A_I1428 (.Y(N450), .A(N6911), .B(N6942));
OAI22XL addgen4_A_I1429 (.Y(N449), .A0(N450), .A1(N438), .B0(N448), .B1(N439));
XNOR2X1 addgen4_A_I1430 (.Y(N452), .A(N6912), .B(N6942));
OAI22XL addgen4_A_I1431 (.Y(N451), .A0(N452), .A1(N438), .B0(N450), .B1(N439));
XNOR2X1 addgen4_A_I1432 (.Y(N454), .A(N6913), .B(N6942));
OAI22XL addgen4_A_I1433 (.Y(N453), .A0(N454), .A1(N438), .B0(N452), .B1(N439));
XNOR2X1 addgen4_A_I1434 (.Y(N456), .A(N6914), .B(N6942));
OAI22XL addgen4_A_I1435 (.Y(N455), .A0(N456), .A1(N438), .B0(N454), .B1(N439));
XNOR2X1 addgen4_A_I1436 (.Y(N458), .A(N6915), .B(N6942));
OAI22XL addgen4_A_I1437 (.Y(N457), .A0(N458), .A1(N438), .B0(N456), .B1(N439));
XNOR2X1 addgen4_A_I1438 (.Y(N460), .A(N6916), .B(N6942));
OAI22XL addgen4_A_I1439 (.Y(N459), .A0(N460), .A1(N438), .B0(N458), .B1(N439));
XNOR2X1 addgen4_A_I1440 (.Y(N462), .A(N6917), .B(N6942));
OAI22XL addgen4_A_I1441 (.Y(N461), .A0(N462), .A1(N438), .B0(N460), .B1(N439));
XNOR2X1 addgen4_A_I1442 (.Y(N464), .A(N6918), .B(N6942));
OAI22XL addgen4_A_I1443 (.Y(N463), .A0(N464), .A1(N438), .B0(N462), .B1(N439));
XNOR2X1 addgen4_A_I1444 (.Y(N466), .A(N6919), .B(N6942));
OAI22XL addgen4_A_I1445 (.Y(N465), .A0(N466), .A1(N438), .B0(N464), .B1(N439));
XNOR2X1 addgen4_A_I1446 (.Y(N468), .A(N6920), .B(N6942));
OAI22XL addgen4_A_I1447 (.Y(N467), .A0(N468), .A1(N438), .B0(N466), .B1(N439));
XNOR2X1 addgen4_A_I1448 (.Y(N470), .A(N6921), .B(N6942));
OAI22XL addgen4_A_I1449 (.Y(N469), .A0(N470), .A1(N438), .B0(N468), .B1(N439));
XNOR2X1 addgen4_A_I1450 (.Y(N472), .A(N6922), .B(N6942));
OAI22XL addgen4_A_I1451 (.Y(N471), .A0(N472), .A1(N438), .B0(N470), .B1(N439));
XNOR2X1 addgen4_A_I1452 (.Y(N474), .A(N6923), .B(N6942));
OAI22XL addgen4_A_I1453 (.Y(N473), .A0(N474), .A1(N438), .B0(N472), .B1(N439));
XNOR2X1 addgen4_A_I1454 (.Y(N476), .A(N6924), .B(N6942));
OAI22XL addgen4_A_I1455 (.Y(N475), .A0(N476), .A1(N438), .B0(N474), .B1(N439));
XNOR2X1 addgen4_A_I1456 (.Y(N478), .A(N6925), .B(N6942));
OAI22XL addgen4_A_I1457 (.Y(N477), .A0(N478), .A1(N438), .B0(N476), .B1(N439));
XNOR2X1 addgen4_A_I1458 (.Y(N480), .A(N6926), .B(N6942));
OAI22XL addgen4_A_I1459 (.Y(N479), .A0(N480), .A1(N438), .B0(N478), .B1(N439));
XNOR2X1 addgen4_A_I1460 (.Y(N482), .A(N6927), .B(N6942));
OAI22XL addgen4_A_I1461 (.Y(N481), .A0(N482), .A1(N438), .B0(N480), .B1(N439));
XNOR2X1 addgen4_A_I1462 (.Y(N484), .A(N6928), .B(N6942));
OAI22XL addgen4_A_I1463 (.Y(N483), .A0(N484), .A1(N438), .B0(N482), .B1(N439));
XNOR2X1 addgen4_A_I1464 (.Y(N486), .A(N6929), .B(N6942));
OAI22XL addgen4_A_I1465 (.Y(N485), .A0(N486), .A1(N438), .B0(N484), .B1(N439));
XNOR2X1 addgen4_A_I1466 (.Y(N488), .A(N6930), .B(N6942));
OAI22XL addgen4_A_I1467 (.Y(N487), .A0(N488), .A1(N438), .B0(N486), .B1(N439));
XNOR2X1 addgen4_A_I1468 (.Y(N490), .A(N6931), .B(N6942));
OAI22XL addgen4_A_I1469 (.Y(N489), .A0(N490), .A1(N438), .B0(N488), .B1(N439));
INVXL addgen4_A_I1470 (.Y(N492), .A(N6942));
OAI22XL addgen4_A_I1471 (.Y(N491), .A0(N492), .A1(N438), .B0(N490), .B1(N439));
MXI2XL inst_cellmath__24_0_I145 (.Y(N493), .A(N439), .B(N438), .S0(N492));
AOI21XL inst_cellmath__24_0_I146 (.Y(N497), .A0(N438), .A1(N439), .B0(N6942));
XNOR2X1 enc3_A_I1472 (.Y(N502), .A(inst_cellmath__24_0_in0[4]), .B(inst_cellmath__24_0_in0[3]));
XOR2XL enc3_A_I1473 (.Y(N2964), .A(inst_cellmath__24_0_in0[5]), .B(inst_cellmath__24_0_in0[3]));
NAND2X1 enc3_A_I1475 (.Y(N503), .A(N2964), .B(N502));
INVXL inst_cellmath__24_0_I2296 (.Y(N6947), .A(inst_cellmath__24_0_in0[5]));
NAND2XL inst_cellmath__24_0_I151 (.Y(N507), .A(inst_cellmath__24_0_in0[3]), .B(inst_cellmath__24_0_in0[4]));
AND2XL inst_cellmath__24_0_I152 (.Y(N508), .A(inst_cellmath__24_0_in0[5]), .B(N507));
XNOR2X1 addgen4_A_I1476 (.Y(N510), .A(N6909), .B(N6947));
OAI22XL addgen4_A_I1477 (.Y(N509), .A0(N510), .A1(N502), .B0(N6947), .B1(N503));
XNOR2X1 addgen4_A_I1478 (.Y(N512), .A(N6910), .B(N6947));
OAI22XL addgen4_A_I1479 (.Y(N511), .A0(N512), .A1(N502), .B0(N510), .B1(N503));
XNOR2X1 addgen4_A_I1480 (.Y(N514), .A(N6911), .B(N6947));
OAI22XL addgen4_A_I1481 (.Y(N513), .A0(N514), .A1(N502), .B0(N512), .B1(N503));
XNOR2X1 addgen4_A_I1482 (.Y(N516), .A(N6912), .B(N6947));
OAI22XL addgen4_A_I1483 (.Y(N515), .A0(N516), .A1(N502), .B0(N514), .B1(N503));
XNOR2X1 addgen4_A_I1484 (.Y(N518), .A(N6913), .B(N6947));
OAI22XL addgen4_A_I1485 (.Y(N517), .A0(N518), .A1(N502), .B0(N516), .B1(N503));
XNOR2X1 addgen4_A_I1486 (.Y(N520), .A(N6914), .B(N6947));
OAI22XL addgen4_A_I1487 (.Y(N519), .A0(N520), .A1(N502), .B0(N518), .B1(N503));
XNOR2X1 addgen4_A_I1488 (.Y(N522), .A(N6915), .B(N6947));
OAI22XL addgen4_A_I1489 (.Y(N521), .A0(N522), .A1(N502), .B0(N520), .B1(N503));
XNOR2X1 addgen4_A_I1490 (.Y(N524), .A(N6916), .B(N6947));
OAI22XL addgen4_A_I1491 (.Y(N523), .A0(N524), .A1(N502), .B0(N522), .B1(N503));
XNOR2X1 addgen4_A_I1492 (.Y(N526), .A(N6917), .B(N6947));
OAI22XL addgen4_A_I1493 (.Y(N525), .A0(N526), .A1(N502), .B0(N524), .B1(N503));
XNOR2X1 addgen4_A_I1494 (.Y(N528), .A(N6918), .B(N6947));
OAI22XL addgen4_A_I1495 (.Y(N527), .A0(N528), .A1(N502), .B0(N526), .B1(N503));
XNOR2X1 addgen4_A_I1496 (.Y(N530), .A(N6919), .B(N6947));
OAI22XL addgen4_A_I1497 (.Y(N529), .A0(N530), .A1(N502), .B0(N528), .B1(N503));
XNOR2X1 addgen4_A_I1498 (.Y(N532), .A(N6920), .B(N6947));
OAI22XL addgen4_A_I1499 (.Y(N531), .A0(N532), .A1(N502), .B0(N530), .B1(N503));
XNOR2X1 addgen4_A_I1500 (.Y(N534), .A(N6921), .B(N6947));
OAI22XL addgen4_A_I1501 (.Y(N533), .A0(N534), .A1(N502), .B0(N532), .B1(N503));
XNOR2X1 addgen4_A_I1502 (.Y(N536), .A(N6922), .B(N6947));
OAI22XL addgen4_A_I1503 (.Y(N535), .A0(N536), .A1(N502), .B0(N534), .B1(N503));
XNOR2X1 addgen4_A_I1504 (.Y(N538), .A(N6923), .B(N6947));
OAI22XL addgen4_A_I1505 (.Y(N537), .A0(N538), .A1(N502), .B0(N536), .B1(N503));
XNOR2X1 addgen4_A_I1506 (.Y(N540), .A(N6924), .B(N6947));
OAI22XL addgen4_A_I1507 (.Y(N539), .A0(N540), .A1(N502), .B0(N538), .B1(N503));
XNOR2X1 addgen4_A_I1508 (.Y(N542), .A(N6925), .B(N6947));
OAI22XL addgen4_A_I1509 (.Y(N541), .A0(N542), .A1(N502), .B0(N540), .B1(N503));
XNOR2X1 addgen4_A_I1510 (.Y(N544), .A(N6926), .B(N6947));
OAI22XL addgen4_A_I1511 (.Y(N543), .A0(N544), .A1(N502), .B0(N542), .B1(N503));
XNOR2X1 addgen4_A_I1512 (.Y(N546), .A(N6927), .B(N6947));
OAI22XL addgen4_A_I1513 (.Y(N545), .A0(N546), .A1(N502), .B0(N544), .B1(N503));
XNOR2X1 addgen4_A_I1514 (.Y(N548), .A(N6928), .B(N6947));
OAI22XL addgen4_A_I1515 (.Y(N547), .A0(N548), .A1(N502), .B0(N546), .B1(N503));
XNOR2X1 addgen4_A_I1516 (.Y(N550), .A(N6929), .B(N6947));
OAI22XL addgen4_A_I1517 (.Y(N549), .A0(N550), .A1(N502), .B0(N548), .B1(N503));
XNOR2X1 addgen4_A_I1518 (.Y(N552), .A(N6930), .B(N6947));
OAI22XL addgen4_A_I1519 (.Y(N551), .A0(N552), .A1(N502), .B0(N550), .B1(N503));
XNOR2X1 addgen4_A_I1520 (.Y(N554), .A(N6931), .B(N6947));
OAI22XL addgen4_A_I1521 (.Y(N553), .A0(N554), .A1(N502), .B0(N552), .B1(N503));
INVXL addgen4_A_I1522 (.Y(N556), .A(N6947));
OAI22XL addgen4_A_I1523 (.Y(N555), .A0(N556), .A1(N502), .B0(N554), .B1(N503));
MXI2XL inst_cellmath__24_0_I177 (.Y(N557), .A(N503), .B(N502), .S0(N556));
AOI21XL inst_cellmath__24_0_I178 (.Y(N561), .A0(N502), .A1(N503), .B0(N6947));
XNOR2X1 enc3_A_I1524 (.Y(N566), .A(inst_cellmath__24_0_in0[6]), .B(inst_cellmath__24_0_in0[5]));
XOR2XL enc3_A_I1525 (.Y(N3191), .A(inst_cellmath__24_0_in0[7]), .B(inst_cellmath__24_0_in0[5]));
NAND2X1 enc3_A_I1527 (.Y(N567), .A(N3191), .B(N566));
INVXL inst_cellmath__24_0_I2301 (.Y(N6952), .A(inst_cellmath__24_0_in0[7]));
NAND2XL inst_cellmath__24_0_I183 (.Y(N571), .A(inst_cellmath__24_0_in0[5]), .B(inst_cellmath__24_0_in0[6]));
AND2XL inst_cellmath__24_0_I184 (.Y(N572), .A(inst_cellmath__24_0_in0[7]), .B(N571));
XNOR2X1 addgen4_A_I1528 (.Y(N574), .A(N6909), .B(N6952));
OAI22XL addgen4_A_I1529 (.Y(N573), .A0(N574), .A1(N566), .B0(N6952), .B1(N567));
XNOR2X1 addgen4_A_I1530 (.Y(N576), .A(N6910), .B(N6952));
OAI22XL addgen4_A_I1531 (.Y(N575), .A0(N576), .A1(N566), .B0(N574), .B1(N567));
XNOR2X1 addgen4_A_I1532 (.Y(N578), .A(N6911), .B(N6952));
OAI22XL addgen4_A_I1533 (.Y(N577), .A0(N578), .A1(N566), .B0(N576), .B1(N567));
XNOR2X1 addgen4_A_I1534 (.Y(N580), .A(N6912), .B(N6952));
OAI22XL addgen4_A_I1535 (.Y(N579), .A0(N580), .A1(N566), .B0(N578), .B1(N567));
XNOR2X1 addgen4_A_I1536 (.Y(N582), .A(N6913), .B(N6952));
OAI22XL addgen4_A_I1537 (.Y(N581), .A0(N582), .A1(N566), .B0(N580), .B1(N567));
XNOR2X1 addgen4_A_I1538 (.Y(N584), .A(N6914), .B(N6952));
OAI22XL addgen4_A_I1539 (.Y(N583), .A0(N584), .A1(N566), .B0(N582), .B1(N567));
XNOR2X1 addgen4_A_I1540 (.Y(N586), .A(N6915), .B(N6952));
OAI22XL addgen4_A_I1541 (.Y(N585), .A0(N586), .A1(N566), .B0(N584), .B1(N567));
XNOR2X1 addgen4_A_I1542 (.Y(N588), .A(N6916), .B(N6952));
OAI22XL addgen4_A_I1543 (.Y(N587), .A0(N588), .A1(N566), .B0(N586), .B1(N567));
XNOR2X1 addgen4_A_I1544 (.Y(N590), .A(N6917), .B(N6952));
OAI22XL addgen4_A_I1545 (.Y(N589), .A0(N590), .A1(N566), .B0(N588), .B1(N567));
XNOR2X1 addgen4_A_I1546 (.Y(N592), .A(N6918), .B(N6952));
OAI22XL addgen4_A_I1547 (.Y(N591), .A0(N592), .A1(N566), .B0(N590), .B1(N567));
XNOR2X1 addgen4_A_I1548 (.Y(N594), .A(N6919), .B(N6952));
OAI22XL addgen4_A_I1549 (.Y(N593), .A0(N594), .A1(N566), .B0(N592), .B1(N567));
XNOR2X1 addgen4_A_I1550 (.Y(N596), .A(N6920), .B(N6952));
OAI22XL addgen4_A_I1551 (.Y(N595), .A0(N596), .A1(N566), .B0(N594), .B1(N567));
XNOR2X1 addgen4_A_I1552 (.Y(N598), .A(N6921), .B(N6952));
OAI22XL addgen4_A_I1553 (.Y(N597), .A0(N598), .A1(N566), .B0(N596), .B1(N567));
XNOR2X1 addgen4_A_I1554 (.Y(N600), .A(N6922), .B(N6952));
OAI22XL addgen4_A_I1555 (.Y(N599), .A0(N600), .A1(N566), .B0(N598), .B1(N567));
XNOR2X1 addgen4_A_I1556 (.Y(N602), .A(N6923), .B(N6952));
OAI22XL addgen4_A_I1557 (.Y(N601), .A0(N602), .A1(N566), .B0(N600), .B1(N567));
XNOR2X1 addgen4_A_I1558 (.Y(N604), .A(N6924), .B(N6952));
OAI22XL addgen4_A_I1559 (.Y(N603), .A0(N604), .A1(N566), .B0(N602), .B1(N567));
XNOR2X1 addgen4_A_I1560 (.Y(N606), .A(N6925), .B(N6952));
OAI22XL addgen4_A_I1561 (.Y(N605), .A0(N606), .A1(N566), .B0(N604), .B1(N567));
XNOR2X1 addgen4_A_I1562 (.Y(N608), .A(N6926), .B(N6952));
OAI22XL addgen4_A_I1563 (.Y(N607), .A0(N608), .A1(N566), .B0(N606), .B1(N567));
XNOR2X1 addgen4_A_I1564 (.Y(N610), .A(N6927), .B(N6952));
OAI22XL addgen4_A_I1565 (.Y(N609), .A0(N610), .A1(N566), .B0(N608), .B1(N567));
XNOR2X1 addgen4_A_I1566 (.Y(N612), .A(N6928), .B(N6952));
OAI22XL addgen4_A_I1567 (.Y(N611), .A0(N612), .A1(N566), .B0(N610), .B1(N567));
XNOR2X1 addgen4_A_I1568 (.Y(N614), .A(N6929), .B(N6952));
OAI22XL addgen4_A_I1569 (.Y(N613), .A0(N614), .A1(N566), .B0(N612), .B1(N567));
XNOR2X1 addgen4_A_I1570 (.Y(N616), .A(N6930), .B(N6952));
OAI22XL addgen4_A_I1571 (.Y(N615), .A0(N616), .A1(N566), .B0(N614), .B1(N567));
XNOR2X1 addgen4_A_I1572 (.Y(N618), .A(N6931), .B(N6952));
OAI22XL addgen4_A_I1573 (.Y(N617), .A0(N618), .A1(N566), .B0(N616), .B1(N567));
INVXL addgen4_A_I1574 (.Y(N620), .A(N6952));
OAI22XL addgen4_A_I1575 (.Y(N619), .A0(N620), .A1(N566), .B0(N618), .B1(N567));
MXI2XL inst_cellmath__24_0_I209 (.Y(N621), .A(N567), .B(N566), .S0(N620));
AOI21XL inst_cellmath__24_0_I210 (.Y(N625), .A0(N566), .A1(N567), .B0(N6952));
XNOR2X1 enc3_A_I1576 (.Y(N630), .A(inst_cellmath__24_0_in0[8]), .B(inst_cellmath__24_0_in0[7]));
XOR2XL enc3_A_I1577 (.Y(N3418), .A(inst_cellmath__24_0_in0[9]), .B(inst_cellmath__24_0_in0[7]));
NAND2X1 enc3_A_I1579 (.Y(N631), .A(N3418), .B(N630));
INVXL inst_cellmath__24_0_I2306 (.Y(N6957), .A(inst_cellmath__24_0_in0[9]));
NAND2XL inst_cellmath__24_0_I215 (.Y(N635), .A(inst_cellmath__24_0_in0[7]), .B(inst_cellmath__24_0_in0[8]));
AND2XL inst_cellmath__24_0_I216 (.Y(N636), .A(inst_cellmath__24_0_in0[9]), .B(N635));
XNOR2X1 addgen4_A_I1580 (.Y(N638), .A(N6909), .B(N6957));
OAI22XL addgen4_A_I1581 (.Y(N637), .A0(N638), .A1(N630), .B0(N6957), .B1(N631));
XNOR2X1 addgen4_A_I1582 (.Y(N640), .A(N6910), .B(N6957));
OAI22XL addgen4_A_I1583 (.Y(N639), .A0(N640), .A1(N630), .B0(N638), .B1(N631));
XNOR2X1 addgen4_A_I1584 (.Y(N642), .A(N6911), .B(N6957));
OAI22XL addgen4_A_I1585 (.Y(N641), .A0(N642), .A1(N630), .B0(N640), .B1(N631));
XNOR2X1 addgen4_A_I1586 (.Y(N644), .A(N6912), .B(N6957));
OAI22XL addgen4_A_I1587 (.Y(N643), .A0(N644), .A1(N630), .B0(N642), .B1(N631));
XNOR2X1 addgen4_A_I1588 (.Y(N646), .A(N6913), .B(N6957));
OAI22XL addgen4_A_I1589 (.Y(N645), .A0(N646), .A1(N630), .B0(N644), .B1(N631));
XNOR2X1 addgen4_A_I1590 (.Y(N648), .A(N6914), .B(N6957));
OAI22XL addgen4_A_I1591 (.Y(N647), .A0(N648), .A1(N630), .B0(N646), .B1(N631));
XNOR2X1 addgen4_A_I1592 (.Y(N650), .A(N6915), .B(N6957));
OAI22XL addgen4_A_I1593 (.Y(N649), .A0(N650), .A1(N630), .B0(N648), .B1(N631));
XNOR2X1 addgen4_A_I1594 (.Y(N652), .A(N6916), .B(N6957));
OAI22XL addgen4_A_I1595 (.Y(N651), .A0(N652), .A1(N630), .B0(N650), .B1(N631));
XNOR2X1 addgen4_A_I1596 (.Y(N654), .A(N6917), .B(N6957));
OAI22XL addgen4_A_I1597 (.Y(N653), .A0(N654), .A1(N630), .B0(N652), .B1(N631));
XNOR2X1 addgen4_A_I1598 (.Y(N656), .A(N6918), .B(N6957));
OAI22XL addgen4_A_I1599 (.Y(N655), .A0(N656), .A1(N630), .B0(N654), .B1(N631));
XNOR2X1 addgen4_A_I1600 (.Y(N658), .A(N6919), .B(N6957));
OAI22XL addgen4_A_I1601 (.Y(N657), .A0(N658), .A1(N630), .B0(N656), .B1(N631));
XNOR2X1 addgen4_A_I1602 (.Y(N660), .A(N6920), .B(N6957));
OAI22XL addgen4_A_I1603 (.Y(N659), .A0(N660), .A1(N630), .B0(N658), .B1(N631));
XNOR2X1 addgen4_A_I1604 (.Y(N662), .A(N6921), .B(N6957));
OAI22XL addgen4_A_I1605 (.Y(N661), .A0(N662), .A1(N630), .B0(N660), .B1(N631));
XNOR2X1 addgen4_A_I1606 (.Y(N664), .A(N6922), .B(N6957));
OAI22XL addgen4_A_I1607 (.Y(N663), .A0(N664), .A1(N630), .B0(N662), .B1(N631));
XNOR2X1 addgen4_A_I1608 (.Y(N666), .A(N6923), .B(N6957));
OAI22XL addgen4_A_I1609 (.Y(N665), .A0(N666), .A1(N630), .B0(N664), .B1(N631));
XNOR2X1 addgen4_A_I1610 (.Y(N668), .A(N6924), .B(N6957));
OAI22XL addgen4_A_I1611 (.Y(N667), .A0(N668), .A1(N630), .B0(N666), .B1(N631));
XNOR2X1 addgen4_A_I1612 (.Y(N670), .A(N6925), .B(N6957));
OAI22XL addgen4_A_I1613 (.Y(N669), .A0(N670), .A1(N630), .B0(N668), .B1(N631));
XNOR2X1 addgen4_A_I1614 (.Y(N672), .A(N6926), .B(N6957));
OAI22XL addgen4_A_I1615 (.Y(N671), .A0(N672), .A1(N630), .B0(N670), .B1(N631));
XNOR2X1 addgen4_A_I1616 (.Y(N674), .A(N6927), .B(N6957));
OAI22XL addgen4_A_I1617 (.Y(N673), .A0(N674), .A1(N630), .B0(N672), .B1(N631));
XNOR2X1 addgen4_A_I1618 (.Y(N676), .A(N6928), .B(N6957));
OAI22XL addgen4_A_I1619 (.Y(N675), .A0(N676), .A1(N630), .B0(N674), .B1(N631));
XNOR2X1 addgen4_A_I1620 (.Y(N678), .A(N6929), .B(N6957));
OAI22XL addgen4_A_I1621 (.Y(N677), .A0(N678), .A1(N630), .B0(N676), .B1(N631));
XNOR2X1 addgen4_A_I1622 (.Y(N680), .A(N6930), .B(N6957));
OAI22XL addgen4_A_I1623 (.Y(N679), .A0(N680), .A1(N630), .B0(N678), .B1(N631));
XNOR2X1 addgen4_A_I1624 (.Y(N682), .A(N6931), .B(N6957));
OAI22XL addgen4_A_I1625 (.Y(N681), .A0(N682), .A1(N630), .B0(N680), .B1(N631));
INVXL addgen4_A_I1626 (.Y(N684), .A(N6957));
OAI22XL addgen4_A_I1627 (.Y(N683), .A0(N684), .A1(N630), .B0(N682), .B1(N631));
MXI2XL inst_cellmath__24_0_I241 (.Y(N685), .A(N631), .B(N630), .S0(N684));
AOI21XL inst_cellmath__24_0_I242 (.Y(N689), .A0(N630), .A1(N631), .B0(N6957));
XNOR2X1 enc3_A_I1628 (.Y(N694), .A(inst_cellmath__24_0_in0[10]), .B(inst_cellmath__24_0_in0[9]));
XOR2XL enc3_A_I1629 (.Y(N3645), .A(inst_cellmath__24_0_in0[11]), .B(inst_cellmath__24_0_in0[9]));
NAND2X1 enc3_A_I1631 (.Y(N695), .A(N3645), .B(N694));
INVXL inst_cellmath__24_0_I2311 (.Y(N6962), .A(inst_cellmath__24_0_in0[11]));
NAND2XL inst_cellmath__24_0_I247 (.Y(N699), .A(inst_cellmath__24_0_in0[9]), .B(inst_cellmath__24_0_in0[10]));
AND2XL inst_cellmath__24_0_I248 (.Y(N700), .A(inst_cellmath__24_0_in0[11]), .B(N699));
XNOR2X1 addgen4_A_I1632 (.Y(N702), .A(N6909), .B(N6962));
OAI22XL addgen4_A_I1633 (.Y(N701), .A0(N702), .A1(N694), .B0(N6962), .B1(N695));
XNOR2X1 addgen4_A_I1634 (.Y(N704), .A(N6910), .B(N6962));
OAI22XL addgen4_A_I1635 (.Y(N703), .A0(N704), .A1(N694), .B0(N702), .B1(N695));
XNOR2X1 addgen4_A_I1636 (.Y(N706), .A(N6911), .B(N6962));
OAI22XL addgen4_A_I1637 (.Y(N705), .A0(N706), .A1(N694), .B0(N704), .B1(N695));
XNOR2X1 addgen4_A_I1638 (.Y(N708), .A(N6912), .B(N6962));
OAI22XL addgen4_A_I1639 (.Y(N707), .A0(N708), .A1(N694), .B0(N706), .B1(N695));
XNOR2X1 addgen4_A_I1640 (.Y(N710), .A(N6913), .B(N6962));
OAI22XL addgen4_A_I1641 (.Y(N709), .A0(N710), .A1(N694), .B0(N708), .B1(N695));
XNOR2X1 addgen4_A_I1642 (.Y(N712), .A(N6914), .B(N6962));
OAI22XL addgen4_A_I1643 (.Y(N711), .A0(N712), .A1(N694), .B0(N710), .B1(N695));
XNOR2X1 addgen4_A_I1644 (.Y(N714), .A(N6915), .B(N6962));
OAI22XL addgen4_A_I1645 (.Y(N713), .A0(N714), .A1(N694), .B0(N712), .B1(N695));
XNOR2X1 addgen4_A_I1646 (.Y(N716), .A(N6916), .B(N6962));
OAI22XL addgen4_A_I1647 (.Y(N715), .A0(N716), .A1(N694), .B0(N714), .B1(N695));
XNOR2X1 addgen4_A_I1648 (.Y(N718), .A(N6917), .B(N6962));
OAI22XL addgen4_A_I1649 (.Y(N717), .A0(N718), .A1(N694), .B0(N716), .B1(N695));
XNOR2X1 addgen4_A_I1650 (.Y(N720), .A(N6918), .B(N6962));
OAI22XL addgen4_A_I1651 (.Y(N719), .A0(N720), .A1(N694), .B0(N718), .B1(N695));
XNOR2X1 addgen4_A_I1652 (.Y(N722), .A(N6919), .B(N6962));
OAI22XL addgen4_A_I1653 (.Y(N721), .A0(N722), .A1(N694), .B0(N720), .B1(N695));
XNOR2X1 addgen4_A_I1654 (.Y(N724), .A(N6920), .B(N6962));
OAI22XL addgen4_A_I1655 (.Y(N723), .A0(N724), .A1(N694), .B0(N722), .B1(N695));
XNOR2X1 addgen4_A_I1656 (.Y(N726), .A(N6921), .B(N6962));
OAI22XL addgen4_A_I1657 (.Y(N725), .A0(N726), .A1(N694), .B0(N724), .B1(N695));
XNOR2X1 addgen4_A_I1658 (.Y(N728), .A(N6922), .B(N6962));
OAI22XL addgen4_A_I1659 (.Y(N727), .A0(N728), .A1(N694), .B0(N726), .B1(N695));
XNOR2X1 addgen4_A_I1660 (.Y(N730), .A(N6923), .B(N6962));
OAI22XL addgen4_A_I1661 (.Y(N729), .A0(N730), .A1(N694), .B0(N728), .B1(N695));
XNOR2X1 addgen4_A_I1662 (.Y(N732), .A(N6924), .B(N6962));
OAI22XL addgen4_A_I1663 (.Y(N731), .A0(N732), .A1(N694), .B0(N730), .B1(N695));
XNOR2X1 addgen4_A_I1664 (.Y(N734), .A(N6925), .B(N6962));
OAI22XL addgen4_A_I1665 (.Y(N733), .A0(N734), .A1(N694), .B0(N732), .B1(N695));
XNOR2X1 addgen4_A_I1666 (.Y(N736), .A(N6926), .B(N6962));
OAI22XL addgen4_A_I1667 (.Y(N735), .A0(N736), .A1(N694), .B0(N734), .B1(N695));
XNOR2X1 addgen4_A_I1668 (.Y(N738), .A(N6927), .B(N6962));
OAI22XL addgen4_A_I1669 (.Y(N737), .A0(N738), .A1(N694), .B0(N736), .B1(N695));
XNOR2X1 addgen4_A_I1670 (.Y(N740), .A(N6928), .B(N6962));
OAI22XL addgen4_A_I1671 (.Y(N739), .A0(N740), .A1(N694), .B0(N738), .B1(N695));
XNOR2X1 addgen4_A_I1672 (.Y(N742), .A(N6929), .B(N6962));
OAI22XL addgen4_A_I1673 (.Y(N741), .A0(N742), .A1(N694), .B0(N740), .B1(N695));
XNOR2X1 addgen4_A_I1674 (.Y(N744), .A(N6930), .B(N6962));
OAI22XL addgen4_A_I1675 (.Y(N743), .A0(N744), .A1(N694), .B0(N742), .B1(N695));
XNOR2X1 addgen4_A_I1676 (.Y(N746), .A(N6931), .B(N6962));
OAI22XL addgen4_A_I1677 (.Y(N745), .A0(N746), .A1(N694), .B0(N744), .B1(N695));
INVXL addgen4_A_I1678 (.Y(N748), .A(N6962));
OAI22XL addgen4_A_I1679 (.Y(N747), .A0(N748), .A1(N694), .B0(N746), .B1(N695));
MXI2XL inst_cellmath__24_0_I273 (.Y(N749), .A(N695), .B(N694), .S0(N748));
AOI21XL inst_cellmath__24_0_I274 (.Y(N753), .A0(N694), .A1(N695), .B0(N6962));
XNOR2X1 enc3_A_I1680 (.Y(N758), .A(inst_cellmath__24_0_in0[12]), .B(inst_cellmath__24_0_in0[11]));
XOR2XL enc3_A_I1681 (.Y(N3872), .A(inst_cellmath__24_0_in0[13]), .B(inst_cellmath__24_0_in0[11]));
NAND2X1 enc3_A_I1683 (.Y(N759), .A(N3872), .B(N758));
INVXL inst_cellmath__24_0_I2316 (.Y(N6967), .A(inst_cellmath__24_0_in0[13]));
NAND2XL inst_cellmath__24_0_I279 (.Y(N763), .A(inst_cellmath__24_0_in0[11]), .B(inst_cellmath__24_0_in0[12]));
AND2XL inst_cellmath__24_0_I280 (.Y(N764), .A(inst_cellmath__24_0_in0[13]), .B(N763));
XNOR2X1 addgen4_A_I1684 (.Y(N766), .A(N6909), .B(N6967));
OAI22XL addgen4_A_I1685 (.Y(N765), .A0(N766), .A1(N758), .B0(N6967), .B1(N759));
XNOR2X1 addgen4_A_I1686 (.Y(N768), .A(N6910), .B(N6967));
OAI22XL addgen4_A_I1687 (.Y(N767), .A0(N768), .A1(N758), .B0(N766), .B1(N759));
XNOR2X1 addgen4_A_I1688 (.Y(N770), .A(N6911), .B(N6967));
OAI22XL addgen4_A_I1689 (.Y(N769), .A0(N770), .A1(N758), .B0(N768), .B1(N759));
XNOR2X1 addgen4_A_I1690 (.Y(N772), .A(N6912), .B(N6967));
OAI22XL addgen4_A_I1691 (.Y(N771), .A0(N772), .A1(N758), .B0(N770), .B1(N759));
XNOR2X1 addgen4_A_I1692 (.Y(N774), .A(N6913), .B(N6967));
OAI22XL addgen4_A_I1693 (.Y(N773), .A0(N774), .A1(N758), .B0(N772), .B1(N759));
XNOR2X1 addgen4_A_I1694 (.Y(N776), .A(N6914), .B(N6967));
OAI22XL addgen4_A_I1695 (.Y(N775), .A0(N776), .A1(N758), .B0(N774), .B1(N759));
XNOR2X1 addgen4_A_I1696 (.Y(N778), .A(N6915), .B(N6967));
OAI22XL addgen4_A_I1697 (.Y(N777), .A0(N778), .A1(N758), .B0(N776), .B1(N759));
XNOR2X1 addgen4_A_I1698 (.Y(N780), .A(N6916), .B(N6967));
OAI22XL addgen4_A_I1699 (.Y(N779), .A0(N780), .A1(N758), .B0(N778), .B1(N759));
XNOR2X1 addgen4_A_I1700 (.Y(N782), .A(N6917), .B(N6967));
OAI22XL addgen4_A_I1701 (.Y(N781), .A0(N782), .A1(N758), .B0(N780), .B1(N759));
XNOR2X1 addgen4_A_I1702 (.Y(N784), .A(N6918), .B(N6967));
OAI22XL addgen4_A_I1703 (.Y(N783), .A0(N784), .A1(N758), .B0(N782), .B1(N759));
XNOR2X1 addgen4_A_I1704 (.Y(N786), .A(N6919), .B(N6967));
OAI22XL addgen4_A_I1705 (.Y(N785), .A0(N786), .A1(N758), .B0(N784), .B1(N759));
XNOR2X1 addgen4_A_I1706 (.Y(N788), .A(N6920), .B(N6967));
OAI22XL addgen4_A_I1707 (.Y(N787), .A0(N788), .A1(N758), .B0(N786), .B1(N759));
XNOR2X1 addgen4_A_I1708 (.Y(N790), .A(N6921), .B(N6967));
OAI22XL addgen4_A_I1709 (.Y(N789), .A0(N790), .A1(N758), .B0(N788), .B1(N759));
XNOR2X1 addgen4_A_I1710 (.Y(N792), .A(N6922), .B(N6967));
OAI22XL addgen4_A_I1711 (.Y(N791), .A0(N792), .A1(N758), .B0(N790), .B1(N759));
XNOR2X1 addgen4_A_I1712 (.Y(N794), .A(N6923), .B(N6967));
OAI22XL addgen4_A_I1713 (.Y(N793), .A0(N794), .A1(N758), .B0(N792), .B1(N759));
XNOR2X1 addgen4_A_I1714 (.Y(N796), .A(N6924), .B(N6967));
OAI22XL addgen4_A_I1715 (.Y(N795), .A0(N796), .A1(N758), .B0(N794), .B1(N759));
XNOR2X1 addgen4_A_I1716 (.Y(N798), .A(N6925), .B(N6967));
OAI22XL addgen4_A_I1717 (.Y(N797), .A0(N798), .A1(N758), .B0(N796), .B1(N759));
XNOR2X1 addgen4_A_I1718 (.Y(N800), .A(N6926), .B(N6967));
OAI22XL addgen4_A_I1719 (.Y(N799), .A0(N800), .A1(N758), .B0(N798), .B1(N759));
XNOR2X1 addgen4_A_I1720 (.Y(N802), .A(N6927), .B(N6967));
OAI22XL addgen4_A_I1721 (.Y(N801), .A0(N802), .A1(N758), .B0(N800), .B1(N759));
XNOR2X1 addgen4_A_I1722 (.Y(N804), .A(N6928), .B(N6967));
OAI22XL addgen4_A_I1723 (.Y(N803), .A0(N804), .A1(N758), .B0(N802), .B1(N759));
XNOR2X1 addgen4_A_I1724 (.Y(N806), .A(N6929), .B(N6967));
OAI22XL addgen4_A_I1725 (.Y(N805), .A0(N806), .A1(N758), .B0(N804), .B1(N759));
XNOR2X1 addgen4_A_I1726 (.Y(N808), .A(N6930), .B(N6967));
OAI22XL addgen4_A_I1727 (.Y(N807), .A0(N808), .A1(N758), .B0(N806), .B1(N759));
XNOR2X1 addgen4_A_I1728 (.Y(N810), .A(N6931), .B(N6967));
OAI22XL addgen4_A_I1729 (.Y(N809), .A0(N810), .A1(N758), .B0(N808), .B1(N759));
INVXL addgen4_A_I1730 (.Y(N812), .A(N6967));
OAI22XL addgen4_A_I1731 (.Y(N811), .A0(N812), .A1(N758), .B0(N810), .B1(N759));
MXI2XL inst_cellmath__24_0_I305 (.Y(N813), .A(N759), .B(N758), .S0(N812));
AOI21XL inst_cellmath__24_0_I306 (.Y(N817), .A0(N758), .A1(N759), .B0(N6967));
XNOR2X1 enc3_A_I1732 (.Y(N822), .A(inst_cellmath__24_0_in0[14]), .B(inst_cellmath__24_0_in0[13]));
XOR2XL enc3_A_I1733 (.Y(N4099), .A(inst_cellmath__24_0_in0[15]), .B(inst_cellmath__24_0_in0[13]));
NAND2X1 enc3_A_I1735 (.Y(N823), .A(N4099), .B(N822));
INVXL inst_cellmath__24_0_I2321 (.Y(N6972), .A(inst_cellmath__24_0_in0[15]));
NAND2XL inst_cellmath__24_0_I311 (.Y(N827), .A(inst_cellmath__24_0_in0[13]), .B(inst_cellmath__24_0_in0[14]));
AND2XL inst_cellmath__24_0_I312 (.Y(N828), .A(inst_cellmath__24_0_in0[15]), .B(N827));
XNOR2X1 addgen4_A_I1736 (.Y(N830), .A(N6909), .B(N6972));
OAI22XL addgen4_A_I1737 (.Y(N829), .A0(N830), .A1(N822), .B0(N6972), .B1(N823));
XNOR2X1 addgen4_A_I1738 (.Y(N832), .A(N6910), .B(N6972));
OAI22XL addgen4_A_I1739 (.Y(N831), .A0(N832), .A1(N822), .B0(N830), .B1(N823));
XNOR2X1 addgen4_A_I1740 (.Y(N834), .A(N6911), .B(N6972));
OAI22XL addgen4_A_I1741 (.Y(N833), .A0(N834), .A1(N822), .B0(N832), .B1(N823));
XNOR2X1 addgen4_A_I1742 (.Y(N836), .A(N6912), .B(N6972));
OAI22XL addgen4_A_I1743 (.Y(N835), .A0(N836), .A1(N822), .B0(N834), .B1(N823));
XNOR2X1 addgen4_A_I1744 (.Y(N838), .A(N6913), .B(N6972));
OAI22XL addgen4_A_I1745 (.Y(N837), .A0(N838), .A1(N822), .B0(N836), .B1(N823));
XNOR2X1 addgen4_A_I1746 (.Y(N840), .A(N6914), .B(N6972));
OAI22XL addgen4_A_I1747 (.Y(N839), .A0(N840), .A1(N822), .B0(N838), .B1(N823));
XNOR2X1 addgen4_A_I1748 (.Y(N842), .A(N6915), .B(N6972));
OAI22XL addgen4_A_I1749 (.Y(N841), .A0(N842), .A1(N822), .B0(N840), .B1(N823));
XNOR2X1 addgen4_A_I1750 (.Y(N844), .A(N6916), .B(N6972));
OAI22XL addgen4_A_I1751 (.Y(N843), .A0(N844), .A1(N822), .B0(N842), .B1(N823));
XNOR2X1 addgen4_A_I1752 (.Y(N846), .A(N6917), .B(N6972));
OAI22XL addgen4_A_I1753 (.Y(N845), .A0(N846), .A1(N822), .B0(N844), .B1(N823));
XNOR2X1 addgen4_A_I1754 (.Y(N848), .A(N6918), .B(N6972));
OAI22XL addgen4_A_I1755 (.Y(N847), .A0(N848), .A1(N822), .B0(N846), .B1(N823));
XNOR2X1 addgen4_A_I1756 (.Y(N850), .A(N6919), .B(N6972));
OAI22XL addgen4_A_I1757 (.Y(N849), .A0(N850), .A1(N822), .B0(N848), .B1(N823));
XNOR2X1 addgen4_A_I1758 (.Y(N852), .A(N6920), .B(N6972));
OAI22XL addgen4_A_I1759 (.Y(N851), .A0(N852), .A1(N822), .B0(N850), .B1(N823));
XNOR2X1 addgen4_A_I1760 (.Y(N854), .A(N6921), .B(N6972));
OAI22XL addgen4_A_I1761 (.Y(N853), .A0(N854), .A1(N822), .B0(N852), .B1(N823));
XNOR2X1 addgen4_A_I1762 (.Y(N856), .A(N6922), .B(N6972));
OAI22XL addgen4_A_I1763 (.Y(N855), .A0(N856), .A1(N822), .B0(N854), .B1(N823));
XNOR2X1 addgen4_A_I1764 (.Y(N858), .A(N6923), .B(N6972));
OAI22XL addgen4_A_I1765 (.Y(N857), .A0(N858), .A1(N822), .B0(N856), .B1(N823));
XNOR2X1 addgen4_A_I1766 (.Y(N860), .A(N6924), .B(N6972));
OAI22XL addgen4_A_I1767 (.Y(N859), .A0(N860), .A1(N822), .B0(N858), .B1(N823));
XNOR2X1 addgen4_A_I1768 (.Y(N862), .A(N6925), .B(N6972));
OAI22XL addgen4_A_I1769 (.Y(N861), .A0(N862), .A1(N822), .B0(N860), .B1(N823));
XNOR2X1 addgen4_A_I1770 (.Y(N864), .A(N6926), .B(N6972));
OAI22XL addgen4_A_I1771 (.Y(N863), .A0(N864), .A1(N822), .B0(N862), .B1(N823));
XNOR2X1 addgen4_A_I1772 (.Y(N866), .A(N6927), .B(N6972));
OAI22XL addgen4_A_I1773 (.Y(N865), .A0(N866), .A1(N822), .B0(N864), .B1(N823));
XNOR2X1 addgen4_A_I1774 (.Y(N868), .A(N6928), .B(N6972));
OAI22XL addgen4_A_I1775 (.Y(N867), .A0(N868), .A1(N822), .B0(N866), .B1(N823));
XNOR2X1 addgen4_A_I1776 (.Y(N870), .A(N6929), .B(N6972));
OAI22XL addgen4_A_I1777 (.Y(N869), .A0(N870), .A1(N822), .B0(N868), .B1(N823));
XNOR2X1 addgen4_A_I1778 (.Y(N872), .A(N6930), .B(N6972));
OAI22XL addgen4_A_I1779 (.Y(N871), .A0(N872), .A1(N822), .B0(N870), .B1(N823));
XNOR2X1 addgen4_A_I1780 (.Y(N874), .A(N6931), .B(N6972));
OAI22XL addgen4_A_I1781 (.Y(N873), .A0(N874), .A1(N822), .B0(N872), .B1(N823));
INVXL addgen4_A_I1782 (.Y(N876), .A(N6972));
OAI22XL addgen4_A_I1783 (.Y(N875), .A0(N876), .A1(N822), .B0(N874), .B1(N823));
MXI2XL inst_cellmath__24_0_I337 (.Y(N877), .A(N823), .B(N822), .S0(N876));
AOI21XL inst_cellmath__24_0_I338 (.Y(N881), .A0(N822), .A1(N823), .B0(N6972));
XNOR2X1 enc3_A_I1784 (.Y(N886), .A(inst_cellmath__24_0_in0[16]), .B(inst_cellmath__24_0_in0[15]));
XOR2XL enc3_A_I1785 (.Y(N4326), .A(inst_cellmath__24_0_in0[17]), .B(inst_cellmath__24_0_in0[15]));
NAND2X1 enc3_A_I1787 (.Y(N887), .A(N4326), .B(N886));
INVXL inst_cellmath__24_0_I2326 (.Y(N6977), .A(inst_cellmath__24_0_in0[17]));
NAND2XL inst_cellmath__24_0_I343 (.Y(N891), .A(inst_cellmath__24_0_in0[15]), .B(inst_cellmath__24_0_in0[16]));
AND2XL inst_cellmath__24_0_I344 (.Y(N892), .A(inst_cellmath__24_0_in0[17]), .B(N891));
XNOR2X1 addgen4_A_I1788 (.Y(N894), .A(N6909), .B(N6977));
OAI22XL addgen4_A_I1789 (.Y(N893), .A0(N894), .A1(N886), .B0(N6977), .B1(N887));
XNOR2X1 addgen4_A_I1790 (.Y(N896), .A(N6910), .B(N6977));
OAI22XL addgen4_A_I1791 (.Y(N895), .A0(N896), .A1(N886), .B0(N894), .B1(N887));
XNOR2X1 addgen4_A_I1792 (.Y(N898), .A(N6911), .B(N6977));
OAI22XL addgen4_A_I1793 (.Y(N897), .A0(N898), .A1(N886), .B0(N896), .B1(N887));
XNOR2X1 addgen4_A_I1794 (.Y(N900), .A(N6912), .B(N6977));
OAI22XL addgen4_A_I1795 (.Y(N899), .A0(N900), .A1(N886), .B0(N898), .B1(N887));
XNOR2X1 addgen4_A_I1796 (.Y(N902), .A(N6913), .B(N6977));
OAI22XL addgen4_A_I1797 (.Y(N901), .A0(N902), .A1(N886), .B0(N900), .B1(N887));
XNOR2X1 addgen4_A_I1798 (.Y(N904), .A(N6914), .B(N6977));
OAI22XL addgen4_A_I1799 (.Y(N903), .A0(N904), .A1(N886), .B0(N902), .B1(N887));
XNOR2X1 addgen4_A_I1800 (.Y(N906), .A(N6915), .B(N6977));
OAI22XL addgen4_A_I1801 (.Y(N905), .A0(N906), .A1(N886), .B0(N904), .B1(N887));
XNOR2X1 addgen4_A_I1802 (.Y(N908), .A(N6916), .B(N6977));
OAI22XL addgen4_A_I1803 (.Y(N907), .A0(N908), .A1(N886), .B0(N906), .B1(N887));
XNOR2X1 addgen4_A_I1804 (.Y(N910), .A(N6917), .B(N6977));
OAI22XL addgen4_A_I1805 (.Y(N909), .A0(N910), .A1(N886), .B0(N908), .B1(N887));
XNOR2X1 addgen4_A_I1806 (.Y(N912), .A(N6918), .B(N6977));
OAI22XL addgen4_A_I1807 (.Y(N911), .A0(N912), .A1(N886), .B0(N910), .B1(N887));
XNOR2X1 addgen4_A_I1808 (.Y(N914), .A(N6919), .B(N6977));
OAI22XL addgen4_A_I1809 (.Y(N913), .A0(N914), .A1(N886), .B0(N912), .B1(N887));
XNOR2X1 addgen4_A_I1810 (.Y(N916), .A(N6920), .B(N6977));
OAI22XL addgen4_A_I1811 (.Y(N915), .A0(N916), .A1(N886), .B0(N914), .B1(N887));
XNOR2X1 addgen4_A_I1812 (.Y(N918), .A(N6921), .B(N6977));
OAI22XL addgen4_A_I1813 (.Y(N917), .A0(N918), .A1(N886), .B0(N916), .B1(N887));
XNOR2X1 addgen4_A_I1814 (.Y(N920), .A(N6922), .B(N6977));
OAI22XL addgen4_A_I1815 (.Y(N919), .A0(N920), .A1(N886), .B0(N918), .B1(N887));
XNOR2X1 addgen4_A_I1816 (.Y(N922), .A(N6923), .B(N6977));
OAI22XL addgen4_A_I1817 (.Y(N921), .A0(N922), .A1(N886), .B0(N920), .B1(N887));
XNOR2X1 addgen4_A_I1818 (.Y(N924), .A(N6924), .B(N6977));
OAI22XL addgen4_A_I1819 (.Y(N923), .A0(N924), .A1(N886), .B0(N922), .B1(N887));
XNOR2X1 addgen4_A_I1820 (.Y(N926), .A(N6925), .B(N6977));
OAI22XL addgen4_A_I1821 (.Y(N925), .A0(N926), .A1(N886), .B0(N924), .B1(N887));
XNOR2X1 addgen4_A_I1822 (.Y(N928), .A(N6926), .B(N6977));
OAI22XL addgen4_A_I1823 (.Y(N927), .A0(N928), .A1(N886), .B0(N926), .B1(N887));
XNOR2X1 addgen4_A_I1824 (.Y(N930), .A(N6927), .B(N6977));
OAI22XL addgen4_A_I1825 (.Y(N929), .A0(N930), .A1(N886), .B0(N928), .B1(N887));
XNOR2X1 addgen4_A_I1826 (.Y(N932), .A(N6928), .B(N6977));
OAI22XL addgen4_A_I1827 (.Y(N931), .A0(N932), .A1(N886), .B0(N930), .B1(N887));
XNOR2X1 addgen4_A_I1828 (.Y(N934), .A(N6929), .B(N6977));
OAI22XL addgen4_A_I1829 (.Y(N933), .A0(N934), .A1(N886), .B0(N932), .B1(N887));
XNOR2X1 addgen4_A_I1830 (.Y(N936), .A(N6930), .B(N6977));
OAI22XL addgen4_A_I1831 (.Y(N935), .A0(N936), .A1(N886), .B0(N934), .B1(N887));
XNOR2X1 addgen4_A_I1832 (.Y(N938), .A(N6931), .B(N6977));
OAI22XL addgen4_A_I1833 (.Y(N937), .A0(N938), .A1(N886), .B0(N936), .B1(N887));
INVXL addgen4_A_I1834 (.Y(N940), .A(N6977));
OAI22XL addgen4_A_I1835 (.Y(N939), .A0(N940), .A1(N886), .B0(N938), .B1(N887));
MXI2XL inst_cellmath__24_0_I369 (.Y(N941), .A(N887), .B(N886), .S0(N940));
AOI21XL inst_cellmath__24_0_I370 (.Y(N945), .A0(N886), .A1(N887), .B0(N6977));
XNOR2X1 enc3_A_I1836 (.Y(N950), .A(inst_cellmath__24_0_in0[18]), .B(inst_cellmath__24_0_in0[17]));
XOR2XL enc3_A_I1837 (.Y(N4553), .A(inst_cellmath__24_0_in0[19]), .B(inst_cellmath__24_0_in0[17]));
NAND2X1 enc3_A_I1839 (.Y(N951), .A(N4553), .B(N950));
INVXL inst_cellmath__24_0_I2331 (.Y(N6982), .A(inst_cellmath__24_0_in0[19]));
NAND2XL inst_cellmath__24_0_I375 (.Y(N955), .A(inst_cellmath__24_0_in0[17]), .B(inst_cellmath__24_0_in0[18]));
AND2XL inst_cellmath__24_0_I376 (.Y(N956), .A(inst_cellmath__24_0_in0[19]), .B(N955));
XNOR2X1 addgen4_A_I1840 (.Y(N958), .A(N6909), .B(N6982));
OAI22XL addgen4_A_I1841 (.Y(N957), .A0(N958), .A1(N950), .B0(N6982), .B1(N951));
XNOR2X1 addgen4_A_I1842 (.Y(N960), .A(N6910), .B(N6982));
OAI22XL addgen4_A_I1843 (.Y(N959), .A0(N960), .A1(N950), .B0(N958), .B1(N951));
XNOR2X1 addgen4_A_I1844 (.Y(N962), .A(N6911), .B(N6982));
OAI22XL addgen4_A_I1845 (.Y(N961), .A0(N962), .A1(N950), .B0(N960), .B1(N951));
XNOR2X1 addgen4_A_I1846 (.Y(N964), .A(N6912), .B(N6982));
OAI22XL addgen4_A_I1847 (.Y(N963), .A0(N964), .A1(N950), .B0(N962), .B1(N951));
XNOR2X1 addgen4_A_I1848 (.Y(N966), .A(N6913), .B(N6982));
OAI22XL addgen4_A_I1849 (.Y(N965), .A0(N966), .A1(N950), .B0(N964), .B1(N951));
XNOR2X1 addgen4_A_I1850 (.Y(N968), .A(N6914), .B(N6982));
OAI22XL addgen4_A_I1851 (.Y(N967), .A0(N968), .A1(N950), .B0(N966), .B1(N951));
XNOR2X1 addgen4_A_I1852 (.Y(N970), .A(N6915), .B(N6982));
OAI22XL addgen4_A_I1853 (.Y(N969), .A0(N970), .A1(N950), .B0(N968), .B1(N951));
XNOR2X1 addgen4_A_I1854 (.Y(N972), .A(N6916), .B(N6982));
OAI22XL addgen4_A_I1855 (.Y(N971), .A0(N972), .A1(N950), .B0(N970), .B1(N951));
XNOR2X1 addgen4_A_I1856 (.Y(N974), .A(N6917), .B(N6982));
OAI22XL addgen4_A_I1857 (.Y(N973), .A0(N974), .A1(N950), .B0(N972), .B1(N951));
XNOR2X1 addgen4_A_I1858 (.Y(N976), .A(N6918), .B(N6982));
OAI22XL addgen4_A_I1859 (.Y(N975), .A0(N976), .A1(N950), .B0(N974), .B1(N951));
XNOR2X1 addgen4_A_I1860 (.Y(N978), .A(N6919), .B(N6982));
OAI22XL addgen4_A_I1861 (.Y(N977), .A0(N978), .A1(N950), .B0(N976), .B1(N951));
XNOR2X1 addgen4_A_I1862 (.Y(N980), .A(N6920), .B(N6982));
OAI22XL addgen4_A_I1863 (.Y(N979), .A0(N980), .A1(N950), .B0(N978), .B1(N951));
XNOR2X1 addgen4_A_I1864 (.Y(N982), .A(N6921), .B(N6982));
OAI22XL addgen4_A_I1865 (.Y(N981), .A0(N982), .A1(N950), .B0(N980), .B1(N951));
XNOR2X1 addgen4_A_I1866 (.Y(N984), .A(N6922), .B(N6982));
OAI22XL addgen4_A_I1867 (.Y(N983), .A0(N984), .A1(N950), .B0(N982), .B1(N951));
XNOR2X1 addgen4_A_I1868 (.Y(N986), .A(N6923), .B(N6982));
OAI22XL addgen4_A_I1869 (.Y(N985), .A0(N986), .A1(N950), .B0(N984), .B1(N951));
XNOR2X1 addgen4_A_I1870 (.Y(N988), .A(N6924), .B(N6982));
OAI22XL addgen4_A_I1871 (.Y(N987), .A0(N988), .A1(N950), .B0(N986), .B1(N951));
XNOR2X1 addgen4_A_I1872 (.Y(N990), .A(N6925), .B(N6982));
OAI22XL addgen4_A_I1873 (.Y(N989), .A0(N990), .A1(N950), .B0(N988), .B1(N951));
XNOR2X1 addgen4_A_I1874 (.Y(N992), .A(N6926), .B(N6982));
OAI22XL addgen4_A_I1875 (.Y(N991), .A0(N992), .A1(N950), .B0(N990), .B1(N951));
XNOR2X1 addgen4_A_I1876 (.Y(N994), .A(N6927), .B(N6982));
OAI22XL addgen4_A_I1877 (.Y(N993), .A0(N994), .A1(N950), .B0(N992), .B1(N951));
XNOR2X1 addgen4_A_I1878 (.Y(N996), .A(N6928), .B(N6982));
OAI22XL addgen4_A_I1879 (.Y(N995), .A0(N996), .A1(N950), .B0(N994), .B1(N951));
XNOR2X1 addgen4_A_I1880 (.Y(N998), .A(N6929), .B(N6982));
OAI22XL addgen4_A_I1881 (.Y(N997), .A0(N998), .A1(N950), .B0(N996), .B1(N951));
XNOR2X1 addgen4_A_I1882 (.Y(N1000), .A(N6930), .B(N6982));
OAI22XL addgen4_A_I1883 (.Y(N999), .A0(N1000), .A1(N950), .B0(N998), .B1(N951));
XNOR2X1 addgen4_A_I1884 (.Y(N1002), .A(N6931), .B(N6982));
OAI22XL addgen4_A_I1885 (.Y(N1001), .A0(N1002), .A1(N950), .B0(N1000), .B1(N951));
INVXL addgen4_A_I1886 (.Y(N1004), .A(N6982));
OAI22XL addgen4_A_I1887 (.Y(N1003), .A0(N1004), .A1(N950), .B0(N1002), .B1(N951));
MXI2XL inst_cellmath__24_0_I401 (.Y(N1005), .A(N951), .B(N950), .S0(N1004));
AOI21XL inst_cellmath__24_0_I402 (.Y(N1009), .A0(N950), .A1(N951), .B0(N6982));
XNOR2X1 enc3_A_I1888 (.Y(N1014), .A(inst_cellmath__24_0_in0[20]), .B(inst_cellmath__24_0_in0[19]));
XOR2XL enc3_A_I1889 (.Y(N4780), .A(inst_cellmath__24_0_in0[21]), .B(inst_cellmath__24_0_in0[19]));
NAND2X1 enc3_A_I1891 (.Y(N1015), .A(N4780), .B(N1014));
INVXL inst_cellmath__24_0_I2336 (.Y(N6987), .A(inst_cellmath__24_0_in0[21]));
NAND2XL inst_cellmath__24_0_I407 (.Y(N1019), .A(inst_cellmath__24_0_in0[19]), .B(inst_cellmath__24_0_in0[20]));
AND2XL inst_cellmath__24_0_I408 (.Y(N1020), .A(inst_cellmath__24_0_in0[21]), .B(N1019));
XNOR2X1 addgen4_A_I1892 (.Y(N1022), .A(N6909), .B(N6987));
OAI22XL addgen4_A_I1893 (.Y(N1021), .A0(N1022), .A1(N1014), .B0(N6987), .B1(N1015));
XNOR2X1 addgen4_A_I1894 (.Y(N1024), .A(N6910), .B(N6987));
OAI22XL addgen4_A_I1895 (.Y(N1023), .A0(N1024), .A1(N1014), .B0(N1022), .B1(N1015));
XNOR2X1 addgen4_A_I1896 (.Y(N1026), .A(N6911), .B(N6987));
OAI22XL addgen4_A_I1897 (.Y(N1025), .A0(N1026), .A1(N1014), .B0(N1024), .B1(N1015));
XNOR2X1 addgen4_A_I1898 (.Y(N1028), .A(N6912), .B(N6987));
OAI22XL addgen4_A_I1899 (.Y(N1027), .A0(N1028), .A1(N1014), .B0(N1026), .B1(N1015));
XNOR2X1 addgen4_A_I1900 (.Y(N1030), .A(N6913), .B(N6987));
OAI22XL addgen4_A_I1901 (.Y(N1029), .A0(N1030), .A1(N1014), .B0(N1028), .B1(N1015));
XNOR2X1 addgen4_A_I1902 (.Y(N1032), .A(N6914), .B(N6987));
OAI22XL addgen4_A_I1903 (.Y(N1031), .A0(N1032), .A1(N1014), .B0(N1030), .B1(N1015));
XNOR2X1 addgen4_A_I1904 (.Y(N1034), .A(N6915), .B(N6987));
OAI22XL addgen4_A_I1905 (.Y(N1033), .A0(N1034), .A1(N1014), .B0(N1032), .B1(N1015));
XNOR2X1 addgen4_A_I1906 (.Y(N1036), .A(N6916), .B(N6987));
OAI22XL addgen4_A_I1907 (.Y(N1035), .A0(N1036), .A1(N1014), .B0(N1034), .B1(N1015));
XNOR2X1 addgen4_A_I1908 (.Y(N1038), .A(N6917), .B(N6987));
OAI22XL addgen4_A_I1909 (.Y(N1037), .A0(N1038), .A1(N1014), .B0(N1036), .B1(N1015));
XNOR2X1 addgen4_A_I1910 (.Y(N1040), .A(N6918), .B(N6987));
OAI22XL addgen4_A_I1911 (.Y(N1039), .A0(N1040), .A1(N1014), .B0(N1038), .B1(N1015));
XNOR2X1 addgen4_A_I1912 (.Y(N1042), .A(N6919), .B(N6987));
OAI22XL addgen4_A_I1913 (.Y(N1041), .A0(N1042), .A1(N1014), .B0(N1040), .B1(N1015));
XNOR2X1 addgen4_A_I1914 (.Y(N1044), .A(N6920), .B(N6987));
OAI22XL addgen4_A_I1915 (.Y(N1043), .A0(N1044), .A1(N1014), .B0(N1042), .B1(N1015));
XNOR2X1 addgen4_A_I1916 (.Y(N1046), .A(N6921), .B(N6987));
OAI22XL addgen4_A_I1917 (.Y(N1045), .A0(N1046), .A1(N1014), .B0(N1044), .B1(N1015));
XNOR2X1 addgen4_A_I1918 (.Y(N1048), .A(N6922), .B(N6987));
OAI22XL addgen4_A_I1919 (.Y(N1047), .A0(N1048), .A1(N1014), .B0(N1046), .B1(N1015));
XNOR2X1 addgen4_A_I1920 (.Y(N1050), .A(N6923), .B(N6987));
OAI22XL addgen4_A_I1921 (.Y(N1049), .A0(N1050), .A1(N1014), .B0(N1048), .B1(N1015));
XNOR2X1 addgen4_A_I1922 (.Y(N1052), .A(N6924), .B(N6987));
OAI22XL addgen4_A_I1923 (.Y(N1051), .A0(N1052), .A1(N1014), .B0(N1050), .B1(N1015));
XNOR2X1 addgen4_A_I1924 (.Y(N1054), .A(N6925), .B(N6987));
OAI22XL addgen4_A_I1925 (.Y(N1053), .A0(N1054), .A1(N1014), .B0(N1052), .B1(N1015));
XNOR2X1 addgen4_A_I1926 (.Y(N1056), .A(N6926), .B(N6987));
OAI22XL addgen4_A_I1927 (.Y(N1055), .A0(N1056), .A1(N1014), .B0(N1054), .B1(N1015));
XNOR2X1 addgen4_A_I1928 (.Y(N1058), .A(N6927), .B(N6987));
OAI22XL addgen4_A_I1929 (.Y(N1057), .A0(N1058), .A1(N1014), .B0(N1056), .B1(N1015));
XNOR2X1 addgen4_A_I1930 (.Y(N1060), .A(N6928), .B(N6987));
OAI22XL addgen4_A_I1931 (.Y(N1059), .A0(N1060), .A1(N1014), .B0(N1058), .B1(N1015));
XNOR2X1 addgen4_A_I1932 (.Y(N1062), .A(N6929), .B(N6987));
OAI22XL addgen4_A_I1933 (.Y(N1061), .A0(N1062), .A1(N1014), .B0(N1060), .B1(N1015));
XNOR2X1 addgen4_A_I1934 (.Y(N1064), .A(N6930), .B(N6987));
OAI22XL addgen4_A_I1935 (.Y(N1063), .A0(N1064), .A1(N1014), .B0(N1062), .B1(N1015));
XNOR2X1 addgen4_A_I1936 (.Y(N1066), .A(N6931), .B(N6987));
OAI22XL addgen4_A_I1937 (.Y(N1065), .A0(N1066), .A1(N1014), .B0(N1064), .B1(N1015));
INVXL addgen4_A_I1938 (.Y(N1068), .A(N6987));
OAI22XL addgen4_A_I1939 (.Y(N1067), .A0(N1068), .A1(N1014), .B0(N1066), .B1(N1015));
MXI2XL inst_cellmath__24_0_I433 (.Y(N1069), .A(N1015), .B(N1014), .S0(N1068));
AOI21XL inst_cellmath__24_0_I434 (.Y(N1073), .A0(N1014), .A1(N1015), .B0(N6987));
XNOR2X1 inst_cellmath__24_0_I1940 (.Y(N1078), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
OR2XL inst_cellmath__24_0_I2511 (.Y(N6990), .A(inst_cellmath__24_0_in0[22]), .B(inst_cellmath__24_0_in0[21]));
NAND2XL inst_cellmath__24_0_I439 (.Y(N1084), .A(inst_cellmath__24_0_in0[21]), .B(inst_cellmath__24_0_in0[22]));
INVXL addgen4_A_I1942 (.Y(N1093), .A(N6909));
OAI21XL addgen4_A_I1943 (.Y(N1092), .A0(N1078), .A1(N1093), .B0(N6990));
INVXL addgen4_A_I1944 (.Y(N1095), .A(N6910));
OAI22XL addgen4_A_I1945 (.Y(N1094), .A0(N1095), .A1(N1078), .B0(N1093), .B1(N6990));
INVXL addgen4_A_I1946 (.Y(N1097), .A(N6911));
OAI22XL addgen4_A_I1947 (.Y(N1096), .A0(N1097), .A1(N1078), .B0(N1095), .B1(N6990));
INVXL addgen4_A_I1948 (.Y(N1099), .A(N6912));
OAI22XL addgen4_A_I1949 (.Y(N1098), .A0(N1099), .A1(N1078), .B0(N1097), .B1(N6990));
INVXL addgen4_A_I1950 (.Y(N1101), .A(N6913));
OAI22XL addgen4_A_I1951 (.Y(N1100), .A0(N1101), .A1(N1078), .B0(N1099), .B1(N6990));
INVXL addgen4_A_I1952 (.Y(N1103), .A(N6914));
OAI22XL addgen4_A_I1953 (.Y(N1102), .A0(N1103), .A1(N1078), .B0(N1101), .B1(N6990));
INVXL addgen4_A_I1954 (.Y(N1105), .A(N6915));
OAI22XL addgen4_A_I1955 (.Y(N1104), .A0(N1105), .A1(N1078), .B0(N1103), .B1(N6990));
INVXL addgen4_A_I1956 (.Y(N1107), .A(N6916));
OAI22XL addgen4_A_I1957 (.Y(N1106), .A0(N1107), .A1(N1078), .B0(N1105), .B1(N6990));
INVXL addgen4_A_I1958 (.Y(N1109), .A(N6917));
OAI22XL addgen4_A_I1959 (.Y(N1108), .A0(N1109), .A1(N1078), .B0(N1107), .B1(N6990));
INVXL addgen4_A_I1960 (.Y(N1111), .A(N6918));
OAI22XL addgen4_A_I1961 (.Y(N1110), .A0(N1111), .A1(N1078), .B0(N1109), .B1(N6990));
INVXL addgen4_A_I1962 (.Y(N1113), .A(N6919));
OAI22XL addgen4_A_I1963 (.Y(N1112), .A0(N1113), .A1(N1078), .B0(N1111), .B1(N6990));
INVXL addgen4_A_I1964 (.Y(N1115), .A(N6920));
OAI22XL addgen4_A_I1965 (.Y(N1114), .A0(N1115), .A1(N1078), .B0(N1113), .B1(N6990));
INVXL addgen4_A_I1966 (.Y(N1117), .A(N6921));
OAI22XL addgen4_A_I1967 (.Y(N1116), .A0(N1117), .A1(N1078), .B0(N1115), .B1(N6990));
INVXL addgen4_A_I1968 (.Y(N1119), .A(N6922));
OAI22XL addgen4_A_I1969 (.Y(N1118), .A0(N1119), .A1(N1078), .B0(N1117), .B1(N6990));
INVXL addgen4_A_I1970 (.Y(N1121), .A(N6923));
OAI22XL addgen4_A_I1971 (.Y(N1120), .A0(N1121), .A1(N1078), .B0(N1119), .B1(N6990));
INVXL addgen4_A_I1972 (.Y(N1123), .A(N6924));
OAI22XL addgen4_A_I1973 (.Y(N1122), .A0(N1123), .A1(N1078), .B0(N1121), .B1(N6990));
INVXL addgen4_A_I1974 (.Y(N1125), .A(N6925));
OAI22XL addgen4_A_I1975 (.Y(N1124), .A0(N1125), .A1(N1078), .B0(N1123), .B1(N6990));
INVXL addgen4_A_I1976 (.Y(N1127), .A(N6926));
OAI22XL addgen4_A_I1977 (.Y(N1126), .A0(N1127), .A1(N1078), .B0(N1125), .B1(N6990));
INVXL addgen4_A_I1978 (.Y(N1129), .A(N6927));
OAI22XL addgen4_A_I1979 (.Y(N1128), .A0(N1129), .A1(N1078), .B0(N1127), .B1(N6990));
INVXL addgen4_A_I1980 (.Y(N1131), .A(N6928));
OAI22XL addgen4_A_I1981 (.Y(N1130), .A0(N1131), .A1(N1078), .B0(N1129), .B1(N6990));
INVXL addgen4_A_I1982 (.Y(N1133), .A(N6929));
OAI22XL addgen4_A_I1983 (.Y(N1132), .A0(N1133), .A1(N1078), .B0(N1131), .B1(N6990));
INVXL addgen4_A_I1984 (.Y(N1135), .A(N6930));
OAI22XL addgen4_A_I1985 (.Y(N1134), .A0(N1135), .A1(N1078), .B0(N1133), .B1(N6990));
INVXL addgen4_A_I1986 (.Y(N1137), .A(N6931));
OAI22XL addgen4_A_I1987 (.Y(N1136), .A0(N1137), .A1(N1078), .B0(N1135), .B1(N6990));
NOR2XL inst_cellmath__24_0_I464 (.Y(N1138), .A(N1137), .B(N6990));
INVXL inst_cellmath__24_0_I465 (.Y(N1140), .A(N1078));
NAND2XL inst_cellmath__24_0_I466 (.Y(N1144), .A(N1078), .B(N6990));
INVXL inst_cellmath__24_0_I499 (.Y(N1212), .A(N433));
INVXL inst_cellmath__24_0_I500 (.Y(N1213), .A(N497));
INVXL inst_cellmath__24_0_I501 (.Y(N1214), .A(N561));
INVXL inst_cellmath__24_0_I502 (.Y(N1215), .A(N625));
INVXL inst_cellmath__24_0_I503 (.Y(N1216), .A(N689));
INVXL inst_cellmath__24_0_I504 (.Y(N1217), .A(N753));
INVXL inst_cellmath__24_0_I505 (.Y(N1218), .A(N817));
INVXL inst_cellmath__24_0_I506 (.Y(N1219), .A(N881));
INVXL inst_cellmath__24_0_I507 (.Y(N1220), .A(N945));
INVXL inst_cellmath__24_0_I508 (.Y(N1221), .A(N1009));
INVXL inst_cellmath__24_0_I509 (.Y(N1222), .A(N1073));
ADDHX1 inst_cellmath__24_0_I510 (.CO(N1224), .S(N1223), .A(N444), .B(N385));
ADDHX1 inst_cellmath__24_0_I511 (.CO(N1226), .S(N1225), .A(N387), .B(N447));
ADDHX1 inst_cellmath__24_0_I512 (.CO(N1228), .S(N1227), .A(N508), .B(N389));
ADDFX1 inst_cellmath__24_0_I513 (.CO(N1230), .S(N1229), .A(N509), .B(N449), .CI(N1226));
ADDHX1 inst_cellmath__24_0_I514 (.CO(N1232), .S(N1231), .A(N391), .B(N451));
ADDFX1 inst_cellmath__24_0_I515 (.CO(N1234), .S(N1233), .A(N1228), .B(N511), .CI(N1231));
ADDHX1 inst_cellmath__24_0_I516 (.CO(N1236), .S(N1235), .A(N572), .B(N393));
ADDFX1 arith_dfa_A_I1988 (.CO(N1239), .S(N5216), .A(N513), .B(N453), .CI(N573));
ADDFX1 arith_dfa_A_I1989 (.CO(N1238), .S(N1237), .A(N1232), .B(N1235), .CI(N5216));
ADDHX1 inst_cellmath__24_0_I518 (.CO(N1241), .S(N1240), .A(N395), .B(N455));
ADDFX1 arith_dfa_A_I1990 (.CO(N1244), .S(N5229), .A(N575), .B(N515), .CI(N1236));
ADDFX1 arith_dfa_A_I1991 (.CO(N1243), .S(N1242), .A(N1240), .B(N1239), .CI(N5229));
ADDHX1 inst_cellmath__24_0_I520 (.CO(N1246), .S(N1245), .A(N636), .B(N397));
ADDFX1 inst_cellmath__24_0_I521 (.CO(N1248), .S(N1247), .A(N517), .B(N457), .CI(N577));
ADDFX1 arith_dfa_A_I1992 (.CO(N1251), .S(N5242), .A(N1241), .B(N637), .CI(N1245));
ADDFX1 arith_dfa_A_I1993 (.CO(N1250), .S(N1249), .A(N1244), .B(N1247), .CI(N5242));
ADDHX1 inst_cellmath__24_0_I523 (.CO(N1253), .S(N1252), .A(N399), .B(N459));
ADDFX1 inst_cellmath__24_0_I524 (.CO(N1255), .S(N1254), .A(N579), .B(N519), .CI(N639));
ADDFX1 arith_dfa_A_I1994 (.CO(N1258), .S(N5255), .A(N1252), .B(N1246), .CI(N1248));
ADDFX1 arith_dfa_A_I1995 (.CO(N1257), .S(N1256), .A(N1251), .B(N1254), .CI(N5255));
ADDHX1 inst_cellmath__24_0_I526 (.CO(N1260), .S(N1259), .A(N700), .B(N401));
ADDFX1 arith_dfa_A_I1996 (.CO(N1263), .S(N5268), .A(N521), .B(N461), .CI(N581));
ADDFX1 arith_dfa_A_I1997 (.CO(N1262), .S(N1261), .A(N1259), .B(N1255), .CI(N5268));
ADDFX1 arith_dfa_A_I1998 (.CO(N1266), .S(N5281), .A(N701), .B(N641), .CI(N1253));
ADDFX1 arith_dfa_A_I1999 (.CO(N1265), .S(N1264), .A(N1261), .B(N1258), .CI(N5281));
ADDHX1 inst_cellmath__24_0_I529 (.CO(N1268), .S(N1267), .A(N403), .B(N463));
ADDFX1 arith_dfa_A_I2000 (.CO(N1271), .S(N5294), .A(N583), .B(N523), .CI(N643));
ADDFX1 arith_dfa_A_I2001 (.CO(N1270), .S(N1269), .A(N1267), .B(N1263), .CI(N5294));
ADDFX1 arith_dfa_A_I2002 (.CO(N1274), .S(N5307), .A(N1260), .B(N703), .CI(N1266));
ADDFX1 arith_dfa_A_I2003 (.CO(N1273), .S(N1272), .A(N1269), .B(N1262), .CI(N5307));
ADDHX1 inst_cellmath__24_0_I532 (.CO(N1276), .S(N1275), .A(N764), .B(N405));
ADDFX1 inst_cellmath__24_0_I533 (.CO(N1278), .S(N1277), .A(N525), .B(N465), .CI(N585));
ADDFX1 arith_dfa_A_I2004 (.CO(N1281), .S(N5320), .A(N705), .B(N645), .CI(N765));
ADDFX1 arith_dfa_A_I2005 (.CO(N1280), .S(N1279), .A(N1275), .B(N1271), .CI(N5320));
ADDFX1 arith_dfa_A_I2006 (.CO(N1284), .S(N5333), .A(N1277), .B(N1268), .CI(N1274));
ADDFX1 arith_dfa_A_I2007 (.CO(N1283), .S(N1282), .A(N1270), .B(N1279), .CI(N5333));
ADDHX1 inst_cellmath__24_0_I536 (.CO(N1286), .S(N1285), .A(N407), .B(N467));
ADDFX1 inst_cellmath__24_0_I537 (.CO(N1288), .S(N1287), .A(N587), .B(N527), .CI(N647));
ADDFX1 arith_dfa_A_I2008 (.CO(N1291), .S(N5346), .A(N767), .B(N707), .CI(N1276));
ADDFX1 arith_dfa_A_I2009 (.CO(N1290), .S(N1289), .A(N1278), .B(N1287), .CI(N5346));
ADDFX1 arith_dfa_A_I2010 (.CO(N1294), .S(N5359), .A(N1281), .B(N1285), .CI(N1280));
ADDFX1 arith_dfa_A_I2011 (.CO(N1293), .S(N1292), .A(N1284), .B(N1289), .CI(N5359));
ADDHX1 inst_cellmath__24_0_I540 (.CO(N1296), .S(N1295), .A(N828), .B(N409));
ADDFX1 arith_dfa_A_I2012 (.CO(N1299), .S(N5372), .A(N529), .B(N469), .CI(N589));
ADDFX1 arith_dfa_A_I2013 (.CO(N1298), .S(N1297), .A(N1295), .B(N1288), .CI(N5372));
ADDFX1 arith_dfa_A_I2014 (.CO(N1302), .S(N5385), .A(N709), .B(N649), .CI(N769));
ADDFX1 arith_dfa_A_I2015 (.CO(N1301), .S(N1300), .A(N829), .B(N1286), .CI(N5385));
ADDFX1 arith_dfa_A_I2016 (.CO(N1305), .S(N5398), .A(N1290), .B(N1291), .CI(N1297));
ADDFX1 arith_dfa_A_I2017 (.CO(N1304), .S(N1303), .A(N1300), .B(N1294), .CI(N5398));
ADDHX1 inst_cellmath__24_0_I544 (.CO(N1307), .S(N1306), .A(N411), .B(N471));
ADDFX1 arith_dfa_A_I2018 (.CO(N1310), .S(N5411), .A(N591), .B(N531), .CI(N651));
ADDFX1 arith_dfa_A_I2019 (.CO(N1309), .S(N1308), .A(N1302), .B(N1299), .CI(N5411));
ADDFX1 arith_dfa_A_I2020 (.CO(N1313), .S(N5424), .A(N771), .B(N711), .CI(N831));
ADDFX1 arith_dfa_A_I2021 (.CO(N1312), .S(N1311), .A(N1296), .B(N1306), .CI(N5424));
ADDFX1 arith_dfa_A_I2022 (.CO(N1316), .S(N5437), .A(N1301), .B(N1298), .CI(N1308));
ADDFX1 arith_dfa_A_I2023 (.CO(N1315), .S(N1314), .A(N1311), .B(N1305), .CI(N5437));
ADDHX1 inst_cellmath__24_0_I548 (.CO(N1318), .S(N1317), .A(N892), .B(N413));
ADDFX1 inst_cellmath__24_0_I549 (.CO(N1320), .S(N1319), .A(N533), .B(N473), .CI(N593));
ADDFX1 arith_dfa_A_I2024 (.CO(N1323), .S(N5450), .A(N713), .B(N653), .CI(N773));
ADDFX1 arith_dfa_A_I2025 (.CO(N1322), .S(N1321), .A(N1313), .B(N1310), .CI(N5450));
ADDFX1 arith_dfa_A_I2026 (.CO(N1326), .S(N5463), .A(N893), .B(N833), .CI(N1307));
ADDFX1 arith_dfa_A_I2027 (.CO(N1325), .S(N1324), .A(N1317), .B(N1319), .CI(N5463));
ADDFX1 arith_dfa_A_I2028 (.CO(N1329), .S(N5476), .A(N1312), .B(N1309), .CI(N1321));
ADDFX1 arith_dfa_A_I2029 (.CO(N1328), .S(N1327), .A(N1324), .B(N1316), .CI(N5476));
ADDHX1 inst_cellmath__24_0_I553 (.CO(N1331), .S(N1330), .A(N415), .B(N475));
ADDFX1 inst_cellmath__24_0_I554 (.CO(N1333), .S(N1332), .A(N595), .B(N535), .CI(N655));
ADDFX1 arith_dfa_A_I2030 (.CO(N1336), .S(N5489), .A(N775), .B(N715), .CI(N835));
ADDFX1 arith_dfa_A_I2031 (.CO(N1335), .S(N1334), .A(N1323), .B(N1320), .CI(N5489));
ADDFX1 arith_dfa_A_I2032 (.CO(N1339), .S(N5502), .A(N1318), .B(N895), .CI(N1330));
ADDFX1 arith_dfa_A_I2033 (.CO(N1338), .S(N1337), .A(N1326), .B(N1332), .CI(N5502));
ADDFX1 arith_dfa_A_I2034 (.CO(N1342), .S(N5515), .A(N1325), .B(N1322), .CI(N1334));
ADDFX1 arith_dfa_A_I2035 (.CO(N1341), .S(N1340), .A(N1337), .B(N1329), .CI(N5515));
ADDHX1 inst_cellmath__24_0_I558 (.CO(N1344), .S(N1343), .A(N956), .B(N417));
ADDFX1 arith_dfa_A_I2036 (.CO(N1347), .S(N5528), .A(N537), .B(N477), .CI(N597));
ADDFX1 arith_dfa_A_I2037 (.CO(N1346), .S(N1345), .A(N1336), .B(N1333), .CI(N5528));
ADDFX1 arith_dfa_A_I2038 (.CO(N1350), .S(N5541), .A(N717), .B(N657), .CI(N777));
ADDFX1 arith_dfa_A_I2039 (.CO(N1349), .S(N1348), .A(N1331), .B(N1343), .CI(N5541));
ADDFX1 arith_dfa_A_I2040 (.CO(N1353), .S(N5554), .A(N897), .B(N837), .CI(N957));
ADDFX1 arith_dfa_A_I2041 (.CO(N1352), .S(N1351), .A(N1335), .B(N1339), .CI(N5554));
ADDFX1 arith_dfa_A_I2042 (.CO(N1356), .S(N5567), .A(N1338), .B(N1345), .CI(N1348));
ADDFX1 arith_dfa_A_I2043 (.CO(N1355), .S(N1354), .A(N1342), .B(N1351), .CI(N5567));
ADDHX1 inst_cellmath__24_0_I563 (.CO(N1358), .S(N1357), .A(N419), .B(N479));
ADDFX1 arith_dfa_A_I2044 (.CO(N1361), .S(N5580), .A(N599), .B(N539), .CI(N659));
ADDFX1 arith_dfa_A_I2045 (.CO(N1360), .S(N1359), .A(N1350), .B(N1347), .CI(N5580));
ADDFX1 arith_dfa_A_I2046 (.CO(N1364), .S(N5593), .A(N779), .B(N719), .CI(N839));
ADDFX1 arith_dfa_A_I2047 (.CO(N1363), .S(N1362), .A(N1357), .B(N1353), .CI(N5593));
ADDFX1 arith_dfa_A_I2048 (.CO(N1367), .S(N5606), .A(N959), .B(N899), .CI(N1344));
ADDFX1 arith_dfa_A_I2049 (.CO(N1366), .S(N1365), .A(N1349), .B(N1346), .CI(N5606));
ADDFX1 arith_dfa_A_I2050 (.CO(N1370), .S(N5619), .A(N1362), .B(N1359), .CI(N1352));
ADDFX1 arith_dfa_A_I2051 (.CO(N1369), .S(N1368), .A(N1365), .B(N1356), .CI(N5619));
ADDHX1 inst_cellmath__24_0_I568 (.CO(N1372), .S(N1371), .A(N1020), .B(N421));
ADDFX1 inst_cellmath__24_0_I569 (.CO(N1374), .S(N1373), .A(N541), .B(N481), .CI(N601));
ADDFX1 arith_dfa_A_I2052 (.CO(N1377), .S(N5632), .A(N721), .B(N661), .CI(N781));
ADDFX1 arith_dfa_A_I2053 (.CO(N1376), .S(N1375), .A(N1364), .B(N1361), .CI(N5632));
ADDFX1 arith_dfa_A_I2054 (.CO(N1380), .S(N5645), .A(N901), .B(N841), .CI(N961));
ADDFX1 arith_dfa_A_I2055 (.CO(N1379), .S(N1378), .A(N1358), .B(N1371), .CI(N5645));
ADDFX1 arith_dfa_A_I2056 (.CO(N1383), .S(N5658), .A(N1367), .B(N1021), .CI(N1373));
ADDFX1 arith_dfa_A_I2057 (.CO(N1382), .S(N1381), .A(N1363), .B(N1360), .CI(N5658));
ADDFX1 arith_dfa_A_I2058 (.CO(N1386), .S(N5671), .A(N1378), .B(N1375), .CI(N1366));
ADDFX1 arith_dfa_A_I2059 (.CO(N1385), .S(N1384), .A(N1370), .B(N1381), .CI(N5671));
ADDHX1 inst_cellmath__24_0_I574 (.CO(N1388), .S(N1387), .A(N423), .B(N483));
ADDFX1 inst_cellmath__24_0_I575 (.CO(N1390), .S(N1389), .A(N603), .B(N543), .CI(N663));
ADDFX1 arith_dfa_A_I2060 (.CO(N1393), .S(N5684), .A(N783), .B(N723), .CI(N843));
ADDFX1 arith_dfa_A_I2061 (.CO(N1392), .S(N1391), .A(N1377), .B(N1374), .CI(N5684));
ADDFX1 arith_dfa_A_I2062 (.CO(N1396), .S(N5697), .A(N963), .B(N903), .CI(N1023));
ADDFX1 arith_dfa_A_I2063 (.CO(N1395), .S(N1394), .A(N1387), .B(N1380), .CI(N5697));
ADDFX1 arith_dfa_A_I2064 (.CO(N1399), .S(N5710), .A(N1389), .B(N1372), .CI(N1376));
ADDFX1 arith_dfa_A_I2065 (.CO(N1398), .S(N1397), .A(N1394), .B(N1391), .CI(N5710));
ADDFX1 arith_dfa_A_I2066 (.CO(N1402), .S(N5723), .A(N1383), .B(N1379), .CI(N1382));
ADDFX1 arith_dfa_A_I2067 (.CO(N1401), .S(N1400), .A(N1386), .B(N1397), .CI(N5723));
ADDHX1 inst_cellmath__24_0_I580 (.CO(N1404), .S(N1403), .A(N1084), .B(N1092));
ADDFX1 arith_dfa_A_I2068 (.CO(N1407), .S(N5736), .A(N425), .B(N1403), .CI(N485));
ADDFX1 arith_dfa_A_I2069 (.CO(N1406), .S(N1405), .A(N1393), .B(N1390), .CI(N5736));
ADDFX1 arith_dfa_A_I2070 (.CO(N1410), .S(N5749), .A(N605), .B(N545), .CI(N665));
ADDFX1 arith_dfa_A_I2071 (.CO(N1409), .S(N1408), .A(N1388), .B(N1396), .CI(N5749));
ADDFX1 arith_dfa_A_I2072 (.CO(N1413), .S(N5762), .A(N785), .B(N725), .CI(N845));
ADDFX1 arith_dfa_A_I2073 (.CO(N1412), .S(N1411), .A(N965), .B(N905), .CI(N5762));
ADDFX1 arith_dfa_A_I2074 (.CO(N1416), .S(N5775), .A(N1392), .B(N1025), .CI(N1395));
ADDFX1 arith_dfa_A_I2075 (.CO(N1415), .S(N1414), .A(N1405), .B(N1399), .CI(N5775));
ADDFX1 arith_dfa_A_I2076 (.CO(N1419), .S(N5788), .A(N1411), .B(N1408), .CI(N1398));
ADDFX1 arith_dfa_A_I2077 (.CO(N1418), .S(N1417), .A(N1402), .B(N1414), .CI(N5788));
ADDHX1 inst_cellmath__24_0_I586 (.CO(N1421), .S(N1420), .A(N1094), .B(N1404));
ADDFX1 arith_dfa_A_I2078 (.CO(N1424), .S(N5801), .A(N427), .B(N1420), .CI(N487));
ADDFX1 arith_dfa_A_I2079 (.CO(N1423), .S(N1422), .A(N1410), .B(N1407), .CI(N5801));
ADDFX1 arith_dfa_A_I2080 (.CO(N1427), .S(N5814), .A(N607), .B(N547), .CI(N667));
ADDFX1 arith_dfa_A_I2081 (.CO(N1426), .S(N1425), .A(N727), .B(N1413), .CI(N5814));
ADDFX1 arith_dfa_A_I2082 (.CO(N1430), .S(N5827), .A(N847), .B(N787), .CI(N907));
ADDFX1 arith_dfa_A_I2083 (.CO(N1429), .S(N1428), .A(N1027), .B(N967), .CI(N5827));
ADDFX1 arith_dfa_A_I2084 (.CO(N1433), .S(N5840), .A(N1409), .B(N1406), .CI(N1412));
ADDFX1 arith_dfa_A_I2085 (.CO(N1432), .S(N1431), .A(N1422), .B(N1416), .CI(N5840));
ADDFX1 arith_dfa_A_I2086 (.CO(N1436), .S(N5853), .A(N1428), .B(N1425), .CI(N1415));
ADDFX1 arith_dfa_A_I2087 (.CO(N1435), .S(N1434), .A(N1431), .B(N1419), .CI(N5853));
ADDFX1 inst_cellmath__24_0_I592 (.CO(N1438), .S(N1437), .A(N1096), .B(N1093), .CI(N1421));
ADDFX1 arith_dfa_A_I2088 (.CO(N1441), .S(N5866), .A(N429), .B(N489), .CI(N549));
ADDFX1 arith_dfa_A_I2089 (.CO(N1440), .S(N1439), .A(N1427), .B(N1424), .CI(N5866));
ADDFX1 arith_dfa_A_I2090 (.CO(N1444), .S(N5879), .A(N669), .B(N609), .CI(N729));
ADDFX1 arith_dfa_A_I2091 (.CO(N1443), .S(N1442), .A(N1437), .B(N1430), .CI(N5879));
ADDFX1 arith_dfa_A_I2092 (.CO(N1447), .S(N5892), .A(N849), .B(N789), .CI(N909));
ADDFX1 arith_dfa_A_I2093 (.CO(N1446), .S(N1445), .A(N1029), .B(N969), .CI(N5892));
ADDFX1 arith_dfa_A_I2094 (.CO(N1450), .S(N5905), .A(N1426), .B(N1423), .CI(N1429));
ADDFX1 arith_dfa_A_I2095 (.CO(N1449), .S(N1448), .A(N1439), .B(N1433), .CI(N5905));
ADDFX1 arith_dfa_A_I2096 (.CO(N1453), .S(N5918), .A(N1445), .B(N1442), .CI(N1432));
ADDFX1 arith_dfa_A_I2097 (.CO(N1452), .S(N1451), .A(N1448), .B(N1436), .CI(N5918));
INVXL fap1_A_I2098 (.Y(N5935), .A(N1095));
ADDFX1 fap1_A_I2099 (.CO(N1455), .S(N1454), .A(N491), .B(N1098), .CI(N5935));
ADDFX1 arith_dfa_A_I2100 (.CO(N1460), .S(N5940), .A(N611), .B(N551), .CI(N671));
ADDFX1 arith_dfa_A_I2101 (.CO(N1459), .S(N1458), .A(N1444), .B(N1441), .CI(N5940));
ADDFX1 arith_dfa_A_I2102 (.CO(N1463), .S(N5953), .A(N791), .B(N731), .CI(N851));
ADDFX1 arith_dfa_A_I2103 (.CO(N1462), .S(N1461), .A(N1438), .B(N1447), .CI(N5953));
ADDFX1 arith_dfa_A_I2104 (.CO(N1466), .S(N5966), .A(N971), .B(N911), .CI(N1031));
ADDFX1 arith_dfa_A_I2105 (.CO(N1465), .S(N1464), .A(N1454), .B(N1212), .CI(N5966));
ADDFX1 arith_dfa_A_I2106 (.CO(N1469), .S(N5979), .A(N1440), .B(N1443), .CI(N1446));
ADDFX1 arith_dfa_A_I2107 (.CO(N1468), .S(N1467), .A(N1464), .B(N1450), .CI(N5979));
ADDFX1 arith_dfa_A_I2108 (.CO(N1472), .S(N5992), .A(N1461), .B(N1458), .CI(N1449));
ADDFX1 arith_dfa_A_I2109 (.CO(N1471), .S(N1470), .A(N1467), .B(N1453), .CI(N5992));
INVXL fap1_A_I2110 (.Y(N6009), .A(N1097));
ADDFX1 fap1_A_I2111 (.CO(N1474), .S(N1473), .A(N1100), .B(N1095), .CI(N6009));
ADDFX1 arith_dfa_A_I2112 (.CO(N1479), .S(N6014), .A(N553), .B(N1473), .CI(N493));
ADDFX1 arith_dfa_A_I2113 (.CO(N1478), .S(N1477), .A(N1460), .B(N1455), .CI(N6014));
ADDFX1 arith_dfa_A_I2114 (.CO(N1482), .S(N6027), .A(N673), .B(N613), .CI(N733));
ADDFX1 arith_dfa_A_I2115 (.CO(N1481), .S(N1480), .A(N1466), .B(N1463), .CI(N6027));
ADDFX1 arith_dfa_A_I2116 (.CO(N1485), .S(N6040), .A(N853), .B(N793), .CI(N913));
ADDFX1 arith_dfa_A_I2117 (.CO(N1484), .S(N1483), .A(N1033), .B(N973), .CI(N6040));
ADDFX1 arith_dfa_A_I2118 (.CO(N1488), .S(N6053), .A(N1465), .B(N1459), .CI(N1462));
ADDFX1 arith_dfa_A_I2119 (.CO(N1487), .S(N1486), .A(N1477), .B(N1469), .CI(N6053));
ADDFX1 arith_dfa_A_I2120 (.CO(N1491), .S(N6066), .A(N1483), .B(N1480), .CI(N1468));
ADDFX1 arith_dfa_A_I2121 (.CO(N1490), .S(N1489), .A(N1486), .B(N1472), .CI(N6066));
ADDFX1 inst_cellmath__24_0_I610 (.CO(N1493), .S(N1492), .A(N1097), .B(N1099), .CI(N1102));
ADDFX1 arith_dfa_A_I2122 (.CO(N1496), .S(N6079), .A(N1492), .B(N1474), .CI(N555));
ADDFX1 arith_dfa_A_I2123 (.CO(N1495), .S(N1494), .A(N615), .B(N1213), .CI(N6079));
ADDFX1 arith_dfa_A_I2124 (.CO(N1499), .S(N6092), .A(N735), .B(N675), .CI(N795));
ADDFX1 arith_dfa_A_I2125 (.CO(N1498), .S(N1497), .A(N1482), .B(N1479), .CI(N6092));
ADDFX1 arith_dfa_A_I2126 (.CO(N1502), .S(N6105), .A(N915), .B(N855), .CI(N975));
ADDFX1 arith_dfa_A_I2127 (.CO(N1501), .S(N1500), .A(N1035), .B(N1485), .CI(N6105));
ADDFX1 arith_dfa_A_I2128 (.CO(N1505), .S(N6118), .A(N1481), .B(N1478), .CI(N1484));
ADDFX1 arith_dfa_A_I2129 (.CO(N1504), .S(N1503), .A(N1497), .B(N1488), .CI(N6118));
ADDFX1 arith_dfa_A_I2130 (.CO(N1508), .S(N6131), .A(N1500), .B(N1494), .CI(N1487));
ADDFX1 arith_dfa_A_I2131 (.CO(N1507), .S(N1506), .A(N1503), .B(N1491), .CI(N6131));
INVXL fap1_A_I2132 (.Y(N6148), .A(N1101));
ADDFX1 fap1_A_I2133 (.CO(N1510), .S(N1509), .A(N1493), .B(N1104), .CI(N6148));
ADDFX1 inst_cellmath__24_0_I617 (.CO(N1514), .S(N1513), .A(N677), .B(N617), .CI(N557));
ADDFX1 arith_dfa_A_I2134 (.CO(N1517), .S(N6153), .A(N797), .B(N737), .CI(N857));
ADDFX1 arith_dfa_A_I2135 (.CO(N1516), .S(N1515), .A(N1502), .B(N1499), .CI(N6153));
ADDFX1 arith_dfa_A_I2136 (.CO(N1520), .S(N6166), .A(N977), .B(N917), .CI(N1037));
ADDFX1 arith_dfa_A_I2137 (.CO(N1519), .S(N1518), .A(N1509), .B(N1496), .CI(N6166));
ADDFX1 arith_dfa_A_I2138 (.CO(N1523), .S(N6179), .A(N1495), .B(N1513), .CI(N1498));
ADDFX1 arith_dfa_A_I2139 (.CO(N1522), .S(N1521), .A(N1515), .B(N1505), .CI(N6179));
ADDFX1 arith_dfa_A_I2140 (.CO(N1526), .S(N6192), .A(N1518), .B(N1501), .CI(N1504));
ADDFX1 arith_dfa_A_I2141 (.CO(N1525), .S(N1524), .A(N1521), .B(N1508), .CI(N6192));
ADDFX1 arith_dfa_A_I2142 (.CO(N1529), .S(N6205), .A(N1101), .B(N1103), .CI(N1106));
ADDFX1 arith_dfa_A_I2143 (.CO(N1528), .S(N1527), .A(N679), .B(N619), .CI(N6205));
ADDFX1 arith_dfa_A_I2144 (.CO(N1532), .S(N6218), .A(N799), .B(N739), .CI(N859));
ADDFX1 arith_dfa_A_I2145 (.CO(N1531), .S(N1530), .A(N1517), .B(N1514), .CI(N6218));
ADDFX1 arith_dfa_A_I2146 (.CO(N1535), .S(N6231), .A(N979), .B(N919), .CI(N1039));
ADDFX1 arith_dfa_A_I2147 (.CO(N1534), .S(N1533), .A(N1214), .B(N1520), .CI(N6231));
ADDFX1 arith_dfa_A_I2148 (.CO(N1538), .S(N6244), .A(N1527), .B(N1510), .CI(N1516));
ADDFX1 arith_dfa_A_I2149 (.CO(N1537), .S(N1536), .A(N1530), .B(N1523), .CI(N6244));
ADDFX1 arith_dfa_A_I2150 (.CO(N1541), .S(N6257), .A(N1533), .B(N1519), .CI(N1522));
ADDFX1 arith_dfa_A_I2151 (.CO(N1540), .S(N1539), .A(N1536), .B(N1526), .CI(N6257));
INVXL fap1_A_I2152 (.Y(N6274), .A(N1105));
ADDFX1 fap1_A_I2153 (.CO(N1543), .S(N1542), .A(N1529), .B(N1108), .CI(N6274));
ADDFX1 arith_dfa_A_I2154 (.CO(N1548), .S(N6279), .A(N621), .B(N681), .CI(N741));
ADDFX1 arith_dfa_A_I2155 (.CO(N1547), .S(N1546), .A(N1532), .B(N1528), .CI(N6279));
ADDFX1 arith_dfa_A_I2156 (.CO(N1551), .S(N6292), .A(N861), .B(N801), .CI(N921));
ADDFX1 arith_dfa_A_I2157 (.CO(N1550), .S(N1549), .A(N1542), .B(N1535), .CI(N6292));
ADDFX1 arith_dfa_A_I2158 (.CO(N1554), .S(N6305), .A(N1041), .B(N981), .CI(N1531));
ADDFX1 arith_dfa_A_I2159 (.CO(N1553), .S(N1552), .A(N1546), .B(N1538), .CI(N6305));
ADDFX1 arith_dfa_A_I2160 (.CO(N1557), .S(N6318), .A(N1549), .B(N1534), .CI(N1537));
ADDFX1 arith_dfa_A_I2161 (.CO(N1556), .S(N1555), .A(N1552), .B(N1541), .CI(N6318));
ADDFX1 inst_cellmath__24_0_I632 (.CO(N1559), .S(N1558), .A(N1105), .B(N1107), .CI(N1110));
ADDFX1 arith_dfa_A_I2162 (.CO(N1562), .S(N6331), .A(N683), .B(N1558), .CI(N743));
ADDFX1 arith_dfa_A_I2163 (.CO(N1561), .S(N1560), .A(N1551), .B(N1548), .CI(N6331));
ADDFX1 arith_dfa_A_I2164 (.CO(N1565), .S(N6344), .A(N863), .B(N803), .CI(N923));
ADDFX1 arith_dfa_A_I2165 (.CO(N1564), .S(N1563), .A(N1543), .B(N1215), .CI(N6344));
ADDFX1 arith_dfa_A_I2166 (.CO(N1568), .S(N6357), .A(N1043), .B(N983), .CI(N1550));
ADDFX1 arith_dfa_A_I2167 (.CO(N1567), .S(N1566), .A(N1560), .B(N1554), .CI(N6357));
ADDFX1 arith_dfa_A_I2168 (.CO(N1571), .S(N6370), .A(N1563), .B(N1547), .CI(N1553));
ADDFX1 arith_dfa_A_I2169 (.CO(N1570), .S(N1569), .A(N1566), .B(N1557), .CI(N6370));
INVXL fap1_A_I2170 (.Y(N6387), .A(N1109));
ADDFX1 fap1_A_I2171 (.CO(N1573), .S(N1572), .A(N1559), .B(N1112), .CI(N6387));
ADDFX1 inst_cellmath__24_0_I638 (.CO(N1577), .S(N1576), .A(N805), .B(N745), .CI(N685));
ADDFX1 arith_dfa_A_I2172 (.CO(N1580), .S(N6392), .A(N925), .B(N865), .CI(N985));
ADDFX1 arith_dfa_A_I2173 (.CO(N1579), .S(N1578), .A(N1565), .B(N1562), .CI(N6392));
ADDFX1 arith_dfa_A_I2174 (.CO(N1583), .S(N6405), .A(N1572), .B(N1045), .CI(N1576));
ADDFX1 arith_dfa_A_I2175 (.CO(N1582), .S(N1581), .A(N1564), .B(N1561), .CI(N6405));
ADDFX1 arith_dfa_A_I2176 (.CO(N1586), .S(N6418), .A(N1568), .B(N1578), .CI(N1581));
ADDFX1 arith_dfa_A_I2177 (.CO(N1585), .S(N1584), .A(N1567), .B(N1571), .CI(N6418));
ADDFX1 arith_dfa_A_I2178 (.CO(N1589), .S(N6431), .A(N1109), .B(N1111), .CI(N1114));
ADDFX1 arith_dfa_A_I2179 (.CO(N1588), .S(N1587), .A(N807), .B(N747), .CI(N6431));
ADDFX1 arith_dfa_A_I2180 (.CO(N1592), .S(N6444), .A(N927), .B(N867), .CI(N987));
ADDFX1 arith_dfa_A_I2181 (.CO(N1591), .S(N1590), .A(N1580), .B(N1577), .CI(N6444));
ADDFX1 arith_dfa_A_I2182 (.CO(N1595), .S(N6457), .A(N1573), .B(N1047), .CI(N1216));
ADDFX1 arith_dfa_A_I2183 (.CO(N1594), .S(N1593), .A(N1579), .B(N1587), .CI(N6457));
ADDFX1 arith_dfa_A_I2184 (.CO(N1598), .S(N6470), .A(N1590), .B(N1583), .CI(N1582));
ADDFX1 arith_dfa_A_I2185 (.CO(N1597), .S(N1596), .A(N1593), .B(N1586), .CI(N6470));
INVXL fap1_A_I2186 (.Y(N6487), .A(N1113));
ADDFX1 fap1_A_I2187 (.CO(N1600), .S(N1599), .A(N1589), .B(N1116), .CI(N6487));
ADDFX1 arith_dfa_A_I2188 (.CO(N1605), .S(N6492), .A(N749), .B(N809), .CI(N869));
ADDFX1 arith_dfa_A_I2189 (.CO(N1604), .S(N1603), .A(N1592), .B(N1588), .CI(N6492));
ADDFX1 arith_dfa_A_I2190 (.CO(N1608), .S(N6505), .A(N989), .B(N929), .CI(N1049));
ADDFX1 arith_dfa_A_I2191 (.CO(N1607), .S(N1606), .A(N1599), .B(N1595), .CI(N6505));
ADDFX1 arith_dfa_A_I2192 (.CO(N1611), .S(N6518), .A(N1606), .B(N1591), .CI(N1603));
ADDFX1 arith_dfa_A_I2193 (.CO(N1610), .S(N1609), .A(N1598), .B(N1594), .CI(N6518));
ADDFX1 inst_cellmath__24_0_I650 (.CO(N1613), .S(N1612), .A(N1113), .B(N1115), .CI(N1118));
ADDFX1 arith_dfa_A_I2194 (.CO(N1616), .S(N6531), .A(N811), .B(N1612), .CI(N871));
ADDFX1 arith_dfa_A_I2195 (.CO(N1615), .S(N1614), .A(N1608), .B(N1605), .CI(N6531));
ADDFX1 arith_dfa_A_I2196 (.CO(N1619), .S(N6544), .A(N991), .B(N931), .CI(N1051));
ADDFX1 arith_dfa_A_I2197 (.CO(N1618), .S(N1617), .A(N1600), .B(N1217), .CI(N6544));
ADDFX1 arith_dfa_A_I2198 (.CO(N1622), .S(N6557), .A(N1604), .B(N1607), .CI(N1614));
ADDFX1 arith_dfa_A_I2199 (.CO(N1621), .S(N1620), .A(N1617), .B(N1611), .CI(N6557));
INVXL fap1_A_I2200 (.Y(N6574), .A(N1117));
ADDFX1 fap1_A_I2201 (.CO(N1624), .S(N1623), .A(N1613), .B(N1120), .CI(N6574));
ADDFX1 inst_cellmath__24_0_I655 (.CO(N1628), .S(N1627), .A(N933), .B(N873), .CI(N813));
ADDFX1 arith_dfa_A_I2202 (.CO(N1631), .S(N6579), .A(N1053), .B(N993), .CI(N1623));
ADDFX1 arith_dfa_A_I2203 (.CO(N1630), .S(N1629), .A(N1616), .B(N1627), .CI(N6579));
ADDFX1 arith_dfa_A_I2204 (.CO(N1634), .S(N6592), .A(N1615), .B(N1619), .CI(N1618));
ADDFX1 arith_dfa_A_I2205 (.CO(N1633), .S(N1632), .A(N1622), .B(N1629), .CI(N6592));
ADDFX1 arith_dfa_A_I2206 (.CO(N1637), .S(N6605), .A(N1117), .B(N1119), .CI(N1122));
ADDFX1 arith_dfa_A_I2207 (.CO(N1636), .S(N1635), .A(N935), .B(N875), .CI(N6605));
ADDFX1 arith_dfa_A_I2208 (.CO(N1640), .S(N6618), .A(N1055), .B(N995), .CI(N1624));
ADDFX1 arith_dfa_A_I2209 (.CO(N1639), .S(N1638), .A(N1218), .B(N1628), .CI(N6618));
ADDFX1 arith_dfa_A_I2210 (.CO(N1643), .S(N6631), .A(N1635), .B(N1631), .CI(N1630));
ADDFX1 arith_dfa_A_I2211 (.CO(N1642), .S(N1641), .A(N1638), .B(N1634), .CI(N6631));
INVXL fap1_A_I2212 (.Y(N6648), .A(N1121));
ADDFX1 fap1_A_I2213 (.CO(N1645), .S(N1644), .A(N1637), .B(N1124), .CI(N6648));
ADDFX1 arith_dfa_A_I2214 (.CO(N1650), .S(N6653), .A(N877), .B(N937), .CI(N997));
ADDFX1 arith_dfa_A_I2215 (.CO(N1649), .S(N1648), .A(N1640), .B(N1636), .CI(N6653));
ADDFX1 arith_dfa_A_I2216 (.CO(N1653), .S(N6666), .A(N1644), .B(N1057), .CI(N1639));
ADDFX1 arith_dfa_A_I2217 (.CO(N1652), .S(N1651), .A(N1648), .B(N1643), .CI(N6666));
ADDFX1 inst_cellmath__24_0_I664 (.CO(N1655), .S(N1654), .A(N1121), .B(N1123), .CI(N1126));
ADDFX1 arith_dfa_A_I2218 (.CO(N1658), .S(N6679), .A(N939), .B(N1654), .CI(N999));
ADDFX1 arith_dfa_A_I2219 (.CO(N1657), .S(N1656), .A(N1219), .B(N1650), .CI(N6679));
ADDFX1 arith_dfa_A_I2220 (.CO(N1661), .S(N6692), .A(N1645), .B(N1059), .CI(N1649));
ADDFX1 arith_dfa_A_I2221 (.CO(N1660), .S(N1659), .A(N1656), .B(N1653), .CI(N6692));
INVXL fap1_A_I2222 (.Y(N6709), .A(N1125));
ADDFX1 fap1_A_I2223 (.CO(N1663), .S(N1662), .A(N1655), .B(N1128), .CI(N6709));
ADDFX1 inst_cellmath__24_0_I668 (.CO(N1667), .S(N1666), .A(N1061), .B(N1001), .CI(N941));
ADDFX1 arith_dfa_A_I2224 (.CO(N1670), .S(N6714), .A(N1658), .B(N1662), .CI(N1666));
ADDFX1 arith_dfa_A_I2225 (.CO(N1669), .S(N1668), .A(N1661), .B(N1657), .CI(N6714));
ADDFX1 arith_dfa_A_I2226 (.CO(N1673), .S(N6727), .A(N1125), .B(N1127), .CI(N1130));
ADDFX1 arith_dfa_A_I2227 (.CO(N1672), .S(N1671), .A(N1063), .B(N1003), .CI(N6727));
ADDFX1 arith_dfa_A_I2228 (.CO(N1676), .S(N6740), .A(N1220), .B(N1663), .CI(N1667));
ADDFX1 arith_dfa_A_I2229 (.CO(N1675), .S(N1674), .A(N1670), .B(N1671), .CI(N6740));
INVXL fap1_A_I2230 (.Y(N6757), .A(N1129));
ADDFX1 fap1_A_I2231 (.CO(N1678), .S(N1677), .A(N1673), .B(N1132), .CI(N6757));
ADDFX1 arith_dfa_A_I2232 (.CO(N1683), .S(N6762), .A(N1005), .B(N1065), .CI(N1677));
ADDFX1 arith_dfa_A_I2233 (.CO(N1682), .S(N1681), .A(N1676), .B(N1672), .CI(N6762));
ADDFX1 inst_cellmath__24_0_I674 (.CO(N1685), .S(N1684), .A(N1129), .B(N1131), .CI(N1134));
ADDFX1 arith_dfa_A_I2234 (.CO(N1688), .S(N6775), .A(N1067), .B(N1684), .CI(N1678));
ADDFX1 arith_dfa_A_I2235 (.CO(N1687), .S(N1686), .A(N1683), .B(N1221), .CI(N6775));
INVXL fap1_A_I2236 (.Y(N6792), .A(N1133));
ADDFX1 fap1_A_I2237 (.CO(N1690), .S(N1689), .A(N1685), .B(N1136), .CI(N6792));
ADDFX1 inst_cellmath__24_0_I677 (.CO(N1694), .S(N1693), .A(N1689), .B(N1069), .CI(N1688));
ADDFX1 arith_dfa_A_I2238 (.CO(N1697), .S(N6797), .A(N1133), .B(N1135), .CI(N1138));
ADDFX1 arith_dfa_A_I2239 (.CO(N1696), .S(N1695), .A(N1222), .B(N1690), .CI(N6797));
ADDFX1 inst_cellmath__24_0_I680 (.CO(N1703), .S(N1702), .A(N1140), .B(N6931), .CI(N1697));
XNOR2X1 inst_cellmath__24_0_I682 (.Y(N1708), .A(N6931), .B(N1144));
NAND2XL inst_cellmath__24_0_I683 (.Y(N1710), .A(inst_cellmath__24_0_in0[1]), .B(N381));
NOR2XL inst_cellmath__24_0_I685 (.Y(N1712), .A(N445), .B(N1223));
NAND2XL inst_cellmath__24_0_I686 (.Y(N1713), .A(N445), .B(N1223));
NOR2XL inst_cellmath__24_0_I687 (.Y(N1714), .A(N1224), .B(N1225));
NAND2XL inst_cellmath__24_0_I688 (.Y(N1715), .A(N1224), .B(N1225));
NOR2XL inst_cellmath__24_0_I689 (.Y(N1716), .A(N1227), .B(N1229));
NAND2XL inst_cellmath__24_0_I690 (.Y(N1717), .A(N1227), .B(N1229));
NOR2XL inst_cellmath__24_0_I691 (.Y(N1718), .A(N1230), .B(N1233));
NAND2XL inst_cellmath__24_0_I692 (.Y(N1719), .A(N1230), .B(N1233));
NOR2XL inst_cellmath__24_0_I693 (.Y(N1720), .A(N1234), .B(N1237));
NAND2XL inst_cellmath__24_0_I694 (.Y(N1721), .A(N1234), .B(N1237));
NOR2XL inst_cellmath__24_0_I695 (.Y(N1722), .A(N1238), .B(N1242));
NAND2XL inst_cellmath__24_0_I696 (.Y(N1723), .A(N1238), .B(N1242));
NOR2XL inst_cellmath__24_0_I697 (.Y(N1724), .A(N1243), .B(N1249));
NAND2XL inst_cellmath__24_0_I698 (.Y(N1725), .A(N1243), .B(N1249));
NOR2XL inst_cellmath__24_0_I699 (.Y(N1726), .A(N1250), .B(N1256));
NAND2XL inst_cellmath__24_0_I700 (.Y(N1727), .A(N1250), .B(N1256));
NOR2XL inst_cellmath__24_0_I701 (.Y(N1728), .A(N1257), .B(N1264));
NAND2XL inst_cellmath__24_0_I702 (.Y(N1729), .A(N1257), .B(N1264));
NOR2XL inst_cellmath__24_0_I703 (.Y(N1730), .A(N1265), .B(N1272));
NAND2XL inst_cellmath__24_0_I704 (.Y(N1731), .A(N1265), .B(N1272));
NOR2XL inst_cellmath__24_0_I705 (.Y(N1732), .A(N1273), .B(N1282));
NAND2XL inst_cellmath__24_0_I706 (.Y(N1733), .A(N1273), .B(N1282));
NOR2XL inst_cellmath__24_0_I707 (.Y(N1734), .A(N1283), .B(N1292));
NAND2XL inst_cellmath__24_0_I708 (.Y(N1735), .A(N1283), .B(N1292));
NOR2XL inst_cellmath__24_0_I709 (.Y(N1736), .A(N1293), .B(N1303));
NAND2XL inst_cellmath__24_0_I710 (.Y(N1737), .A(N1293), .B(N1303));
NOR2XL inst_cellmath__24_0_I711 (.Y(N1738), .A(N1304), .B(N1314));
NAND2XL inst_cellmath__24_0_I712 (.Y(N1739), .A(N1304), .B(N1314));
NOR2XL inst_cellmath__24_0_I713 (.Y(N1740), .A(N1315), .B(N1327));
NAND2XL inst_cellmath__24_0_I714 (.Y(N1741), .A(N1315), .B(N1327));
NOR2XL inst_cellmath__24_0_I715 (.Y(N1742), .A(N1328), .B(N1340));
NAND2XL inst_cellmath__24_0_I716 (.Y(N1743), .A(N1328), .B(N1340));
NOR2XL inst_cellmath__24_0_I717 (.Y(N1744), .A(N1341), .B(N1354));
NAND2XL inst_cellmath__24_0_I718 (.Y(N1745), .A(N1341), .B(N1354));
NOR2XL inst_cellmath__24_0_I721 (.Y(N1748), .A(N6937), .B(N1710));
INVXL inst_cellmath__24_0_I2340 (.Y(N6991), .A(N1712));
INVXL inst_cellmath__24_0_I2341 (.Y(N6992), .A(N1713));
OAI21XL inst_cellmath__24_0_I729 (.Y(N1758), .A0(N6992), .A1(N1748), .B0(N6991));
AOI21XL inst_cellmath__24_0_I737 (.Y(N1766), .A0(N1715), .A1(N1758), .B0(N1714));
INVXL inst_cellmath__24_0_I2348 (.Y(N6999), .A(N1716));
INVXL inst_cellmath__24_0_I2349 (.Y(N7000), .A(N1717));
OAI21XL inst_cellmath__24_0_I749 (.Y(N1778), .A0(N7000), .A1(N1766), .B0(N6999));
AOI21XL inst_cellmath__24_0_I761 (.Y(N1790), .A0(N1719), .A1(N1778), .B0(N1718));
INVXL inst_cellmath__24_0_I2359 (.Y(N7010), .A(N1720));
INVXL inst_cellmath__24_0_I2360 (.Y(N7011), .A(N1721));
OAI21XL inst_cellmath__24_0_I777 (.Y(N1806), .A0(N7011), .A1(N1790), .B0(N7010));
AOI21XL inst_cellmath__24_0_I793 (.Y(N1822), .A0(N1723), .A1(N1806), .B0(N1722));
INVXL inst_cellmath__24_0_I2374 (.Y(N7025), .A(N1724));
INVXL inst_cellmath__24_0_I2375 (.Y(N7026), .A(N1725));
OAI21XL inst_cellmath__24_0_I813 (.Y(N1842), .A0(N7026), .A1(N1822), .B0(N7025));
AOI21XL inst_cellmath__24_0_I833 (.Y(N1862), .A0(N1727), .A1(N1842), .B0(N1726));
AOI21XL inst_cellmath__24_0_I837 (.Y(N1866), .A0(N1731), .A1(N1728), .B0(N1730));
NAND2XL inst_cellmath__24_0_I838 (.Y(N1867), .A(N1731), .B(N1729));
OAI21XL inst_cellmath__24_0_I861 (.Y(N1890), .A0(N1867), .A1(N1862), .B0(N1866));
AO21XL inst_cellmath__24_0_I2512 (.Y(N7064), .A0(N1735), .A1(N1732), .B0(N1734));
AOI21XL inst_cellmath__24_0_I895 (.Y(N1924), .A0(N1733), .A1(N1890), .B0(N1732));
AOI31X1 inst_cellmath__24_0_I2514 (.Y(N1926), .A0(N1735), .A1(N1733), .A2(N1890), .B0(N7064));
AOI21XL inst_cellmath__24_0_I901 (.Y(N1930), .A0(N1739), .A1(N1736), .B0(N1738));
NAND2XL inst_cellmath__24_0_I902 (.Y(N1931), .A(N1739), .B(N1737));
OAI21XL inst_cellmath__24_0_I933 (.Y(N1962), .A0(N1931), .A1(N1926), .B0(N1930));
AOI21XL inst_cellmath__24_0_I937 (.Y(N1966), .A0(N1743), .A1(N1740), .B0(N1742));
NAND2XL inst_cellmath__24_0_I938 (.Y(N1967), .A(N1743), .B(N1741));
INVXL inst_cellmath__24_0_I2449 (.Y(N7100), .A(N1744));
INVXL inst_cellmath__24_0_I2450 (.Y(N7101), .A(N1745));
INVXL inst_cellmath__24_0_I2453 (.Y(N7104), .A(N1966));
INVXL inst_cellmath__24_0_I2454 (.Y(N7105), .A(N1967));
OAI21XL inst_cellmath__24_0_I945 (.Y(N1974), .A0(N7101), .A1(N1966), .B0(N7100));
NOR2XL inst_cellmath__24_0_I946 (.Y(N1975), .A(N7101), .B(N1967));
NOR2BX1 andori2bb1_A_I5136 (.Y(N7162), .AN(N1729), .B(N1862));
NOR2XL andori2bb1_A_I2543 (.Y(N7116), .A(N7162), .B(N1728));
NOR2BX1 andori2bb1_A_I5137 (.Y(N7169), .AN(N1737), .B(N1926));
NOR2XL andori2bb1_A_I2545 (.Y(N7120), .A(N7169), .B(N1736));
AOI21XL inst_cellmath__24_0_I979 (.Y(N2008), .A0(N1741), .A1(N1962), .B0(N1740));
AOI21XL inst_cellmath__24_0_I981 (.Y(N2010), .A0(N7105), .A1(N1962), .B0(N7104));
NAND2BXL inst_cellmath__24_0_I1011 (.Y(N2042), .AN(N1712), .B(N1713));
NAND2BXL inst_cellmath__24_0_I1014 (.Y(N2045), .AN(N1714), .B(N1715));
NAND2BXL inst_cellmath__24_0_I1017 (.Y(N2048), .AN(N1716), .B(N1717));
NAND2BXL inst_cellmath__24_0_I1020 (.Y(N2051), .AN(N1718), .B(N1719));
NAND2BXL inst_cellmath__24_0_I1023 (.Y(N2054), .AN(N1720), .B(N1721));
NAND2BXL inst_cellmath__24_0_I1026 (.Y(N2057), .AN(N1722), .B(N1723));
NAND2BXL inst_cellmath__24_0_I1029 (.Y(N2060), .AN(N1724), .B(N1725));
NAND2BXL inst_cellmath__24_0_I1032 (.Y(N2063), .AN(N1726), .B(N1727));
NAND2BXL inst_cellmath__24_0_I1035 (.Y(N2066), .AN(N1728), .B(N1729));
NAND2BXL inst_cellmath__24_0_I1038 (.Y(N2069), .AN(N1730), .B(N1731));
NAND2BXL inst_cellmath__24_0_I1041 (.Y(N2072), .AN(N1732), .B(N1733));
NAND2BXL inst_cellmath__24_0_I1044 (.Y(N2075), .AN(N1734), .B(N1735));
NAND2BXL inst_cellmath__24_0_I1047 (.Y(N2078), .AN(N1736), .B(N1737));
NAND2BXL inst_cellmath__24_0_I1050 (.Y(N2081), .AN(N1738), .B(N1739));
NAND2BXL inst_cellmath__24_0_I1053 (.Y(N2084), .AN(N1740), .B(N1741));
NAND2BXL inst_cellmath__24_0_I1056 (.Y(N2087), .AN(N1742), .B(N1743));
NAND2BXL inst_cellmath__24_0_I1059 (.Y(N2090), .AN(N1744), .B(N1745));
XOR2XL inst_cellmath__24_0_I1060 (.Y(inst_cellmath__24_0_out0[0]), .A(inst_cellmath__24_0_in0[1]), .B(N381));
XOR2XL inst_cellmath__24_0_I2517 (.Y(inst_cellmath__24_0_out0[1]), .A(N1710), .B(N6937));
XNOR2X1 inst_cellmath__24_0_I1062 (.Y(inst_cellmath__24_0_out0[2]), .A(N1748), .B(N2042));
XOR2XL inst_cellmath__24_0_I2518 (.Y(inst_cellmath__24_0_out0[3]), .A(N1758), .B(N2045));
XNOR2X1 inst_cellmath__24_0_I1064 (.Y(inst_cellmath__24_0_out0[4]), .A(N1766), .B(N2048));
XOR2XL inst_cellmath__24_0_I2519 (.Y(inst_cellmath__24_0_out0[5]), .A(N1778), .B(N2051));
XNOR2X1 inst_cellmath__24_0_I1066 (.Y(inst_cellmath__24_0_out0[6]), .A(N1790), .B(N2054));
XOR2XL inst_cellmath__24_0_I2520 (.Y(inst_cellmath__24_0_out0[7]), .A(N1806), .B(N2057));
XNOR2X1 inst_cellmath__24_0_I1068 (.Y(inst_cellmath__24_0_out0[8]), .A(N1822), .B(N2060));
XOR2XL inst_cellmath__24_0_I2521 (.Y(inst_cellmath__24_0_out0[9]), .A(N1842), .B(N2063));
XNOR2X1 inst_cellmath__24_0_I1070 (.Y(inst_cellmath__24_0_out0[10]), .A(N1862), .B(N2066));
XNOR2X1 inst_cellmath__24_0_I1071 (.Y(inst_cellmath__24_0_out0[11]), .A(N7116), .B(N2069));
XOR2XL inst_cellmath__24_0_I2522 (.Y(inst_cellmath__24_0_out0[12]), .A(N1890), .B(N2072));
XNOR2X1 inst_cellmath__24_0_I1073 (.Y(inst_cellmath__24_0_out0[13]), .A(N1924), .B(N2075));
XNOR2X1 inst_cellmath__24_0_I1074 (.Y(inst_cellmath__24_0_out0[14]), .A(N1926), .B(N2078));
XNOR2X1 inst_cellmath__24_0_I1075 (.Y(inst_cellmath__24_0_out0[15]), .A(N7120), .B(N2081));
XOR2XL inst_cellmath__24_0_I2523 (.Y(inst_cellmath__24_0_out0[16]), .A(N1962), .B(N2084));
XNOR2X1 inst_cellmath__24_0_I1077 (.Y(inst_cellmath__24_0_out0[17]), .A(N2008), .B(N2087));
XNOR2X1 inst_cellmath__24_0_I1078 (.Y(inst_cellmath__24_0_out0[18]), .A(N2010), .B(N2090));
AO21XL inst_cellmath__24_0_I2251 (.Y(N2110), .A0(N1975), .A1(N1962), .B0(N1974));
XOR2XL inst_cellmath__24_0_I1081 (.Y(N2113), .A(N1355), .B(N1368));
NOR2XL inst_cellmath__24_0_I1082 (.Y(N2114), .A(N1369), .B(N1384));
XOR2XL inst_cellmath__24_0_I1083 (.Y(N2115), .A(N1369), .B(N1384));
NOR2XL inst_cellmath__24_0_I1084 (.Y(N2116), .A(N1385), .B(N1400));
XOR2XL inst_cellmath__24_0_I1085 (.Y(N2117), .A(N1385), .B(N1400));
NOR2XL inst_cellmath__24_0_I1086 (.Y(N2118), .A(N1401), .B(N1417));
XOR2XL inst_cellmath__24_0_I1087 (.Y(N2119), .A(N1401), .B(N1417));
NOR2XL inst_cellmath__24_0_I1088 (.Y(N2120), .A(N1418), .B(N1434));
XOR2XL inst_cellmath__24_0_I1089 (.Y(N2121), .A(N1418), .B(N1434));
NOR2XL inst_cellmath__24_0_I1090 (.Y(N2122), .A(N1435), .B(N1451));
XOR2XL inst_cellmath__24_0_I1091 (.Y(N2123), .A(N1435), .B(N1451));
NOR2XL inst_cellmath__24_0_I1092 (.Y(N2124), .A(N1452), .B(N1470));
XOR2XL inst_cellmath__24_0_I1093 (.Y(N2125), .A(N1452), .B(N1470));
NOR2XL inst_cellmath__24_0_I1094 (.Y(N2126), .A(N1471), .B(N1489));
XOR2XL inst_cellmath__24_0_I1095 (.Y(N2127), .A(N1471), .B(N1489));
NOR2XL inst_cellmath__24_0_I1096 (.Y(N2128), .A(N1490), .B(N1506));
XOR2XL inst_cellmath__24_0_I1097 (.Y(N2129), .A(N1490), .B(N1506));
NOR2XL inst_cellmath__24_0_I1098 (.Y(N2130), .A(N1507), .B(N1524));
XOR2XL inst_cellmath__24_0_I1099 (.Y(N2131), .A(N1507), .B(N1524));
NOR2XL inst_cellmath__24_0_I1100 (.Y(N2132), .A(N1525), .B(N1539));
XOR2XL inst_cellmath__24_0_I1101 (.Y(N2133), .A(N1525), .B(N1539));
NOR2XL inst_cellmath__24_0_I1102 (.Y(N2134), .A(N1540), .B(N1555));
XOR2XL inst_cellmath__24_0_I1103 (.Y(N2135), .A(N1540), .B(N1555));
NOR2XL inst_cellmath__24_0_I1104 (.Y(N2136), .A(N1556), .B(N1569));
XOR2XL inst_cellmath__24_0_I1105 (.Y(N2137), .A(N1556), .B(N1569));
NOR2XL inst_cellmath__24_0_I1106 (.Y(N2138), .A(N1570), .B(N1584));
XOR2XL inst_cellmath__24_0_I1107 (.Y(N2139), .A(N1570), .B(N1584));
NOR2XL inst_cellmath__24_0_I1108 (.Y(N2140), .A(N1585), .B(N1596));
XOR2XL inst_cellmath__24_0_I1109 (.Y(N2141), .A(N1585), .B(N1596));
NOR2XL inst_cellmath__24_0_I1110 (.Y(N2142), .A(N1597), .B(N1609));
XOR2XL inst_cellmath__24_0_I1111 (.Y(N2143), .A(N1597), .B(N1609));
NOR2XL inst_cellmath__24_0_I1112 (.Y(N2144), .A(N1620), .B(N1610));
XOR2XL inst_cellmath__24_0_I1113 (.Y(N2145), .A(N1620), .B(N1610));
NOR2XL inst_cellmath__24_0_I1114 (.Y(N2146), .A(N1621), .B(N1632));
XOR2XL inst_cellmath__24_0_I1115 (.Y(N2147), .A(N1621), .B(N1632));
NOR2XL inst_cellmath__24_0_I1116 (.Y(N2148), .A(N1633), .B(N1641));
XOR2XL inst_cellmath__24_0_I1117 (.Y(N2149), .A(N1633), .B(N1641));
NOR2XL inst_cellmath__24_0_I1118 (.Y(N2150), .A(N1642), .B(N1651));
XOR2XL inst_cellmath__24_0_I1119 (.Y(N2151), .A(N1642), .B(N1651));
NOR2XL inst_cellmath__24_0_I1120 (.Y(N2152), .A(N1652), .B(N1659));
XOR2XL inst_cellmath__24_0_I1121 (.Y(N2153), .A(N1652), .B(N1659));
NOR2XL inst_cellmath__24_0_I1122 (.Y(N2154), .A(N1660), .B(N1668));
XOR2XL inst_cellmath__24_0_I1123 (.Y(N2155), .A(N1660), .B(N1668));
NOR2XL inst_cellmath__24_0_I1124 (.Y(N2156), .A(N1674), .B(N1669));
XOR2XL inst_cellmath__24_0_I1125 (.Y(N2157), .A(N1674), .B(N1669));
NOR2XL inst_cellmath__24_0_I1126 (.Y(N2158), .A(N1675), .B(N1681));
XOR2XL inst_cellmath__24_0_I1127 (.Y(N2159), .A(N1675), .B(N1681));
NOR2XL inst_cellmath__24_0_I1128 (.Y(N2160), .A(N1682), .B(N1686));
XOR2XL inst_cellmath__24_0_I1129 (.Y(N2161), .A(N1682), .B(N1686));
NOR2XL inst_cellmath__24_0_I1130 (.Y(N2162), .A(N1693), .B(N1687));
XOR2XL inst_cellmath__24_0_I1131 (.Y(N2163), .A(N1693), .B(N1687));
NOR2XL inst_cellmath__24_0_I1132 (.Y(N2164), .A(N1695), .B(N1694));
XOR2XL inst_cellmath__24_0_I1133 (.Y(N2165), .A(N1695), .B(N1694));
NOR2XL inst_cellmath__24_0_I1134 (.Y(N2166), .A(N1702), .B(N1696));
XOR2XL inst_cellmath__24_0_I1135 (.Y(N2167), .A(N1702), .B(N1696));
XNOR2X1 inst_cellmath__24_0_I1137 (.Y(N2169), .A(N1708), .B(N1703));
AOI2BB2X1 inst_cellmath__24_0_I2252 (.Y(N2170), .A0N(N1355), .A1N(N1368), .B0(N2110), .B1(N2113));
AOI21XL inst_cellmath__24_0_I1140 (.Y(N2172), .A0(N2117), .A1(N2114), .B0(N2116));
NAND2XL inst_cellmath__24_0_I1141 (.Y(N2173), .A(N2117), .B(N2115));
AOI21XL inst_cellmath__24_0_I1142 (.Y(N2174), .A0(N2121), .A1(N2118), .B0(N2120));
NAND2XL inst_cellmath__24_0_I1143 (.Y(N2175), .A(N2121), .B(N2119));
AOI21XL inst_cellmath__24_0_I1144 (.Y(N2176), .A0(N2125), .A1(N2122), .B0(N2124));
NAND2XL inst_cellmath__24_0_I1145 (.Y(N2177), .A(N2125), .B(N2123));
AOI21XL inst_cellmath__24_0_I1146 (.Y(N2178), .A0(N2129), .A1(N2126), .B0(N2128));
NAND2XL inst_cellmath__24_0_I1147 (.Y(N2179), .A(N2129), .B(N2127));
AOI21XL inst_cellmath__24_0_I1148 (.Y(N2180), .A0(N2133), .A1(N2130), .B0(N2132));
NAND2XL inst_cellmath__24_0_I1149 (.Y(N2181), .A(N2133), .B(N2131));
AOI21XL inst_cellmath__24_0_I1150 (.Y(N2182), .A0(N2137), .A1(N2134), .B0(N2136));
NAND2XL inst_cellmath__24_0_I1151 (.Y(N2183), .A(N2137), .B(N2135));
AOI21XL inst_cellmath__24_0_I1152 (.Y(N2184), .A0(N2141), .A1(N2138), .B0(N2140));
NAND2XL inst_cellmath__24_0_I1153 (.Y(N2185), .A(N2141), .B(N2139));
AOI21XL inst_cellmath__24_0_I1154 (.Y(N2186), .A0(N2145), .A1(N2142), .B0(N2144));
NAND2XL inst_cellmath__24_0_I1155 (.Y(N2187), .A(N2145), .B(N2143));
AOI21XL inst_cellmath__24_0_I1156 (.Y(N2188), .A0(N2149), .A1(N2146), .B0(N2148));
NAND2XL inst_cellmath__24_0_I1157 (.Y(N2189), .A(N2149), .B(N2147));
AOI21XL inst_cellmath__24_0_I1158 (.Y(N2190), .A0(N2153), .A1(N2150), .B0(N2152));
NAND2XL inst_cellmath__24_0_I1159 (.Y(N2191), .A(N2153), .B(N2151));
AOI21XL inst_cellmath__24_0_I1160 (.Y(N2192), .A0(N2157), .A1(N2154), .B0(N2156));
NAND2XL inst_cellmath__24_0_I1161 (.Y(N2193), .A(N2157), .B(N2155));
AOI21XL inst_cellmath__24_0_I1162 (.Y(N2194), .A0(N2161), .A1(N2158), .B0(N2160));
NAND2XL inst_cellmath__24_0_I1163 (.Y(N2195), .A(N2161), .B(N2159));
AOI21XL inst_cellmath__24_0_I1164 (.Y(N2196), .A0(N2165), .A1(N2162), .B0(N2164));
NAND2XL inst_cellmath__24_0_I1165 (.Y(N2197), .A(N2165), .B(N2163));
OAI21XL inst_cellmath__24_0_I1168 (.Y(N2200), .A0(N2173), .A1(N2170), .B0(N2172));
OAI21XL inst_cellmath__24_0_I1170 (.Y(N2202), .A0(N2177), .A1(N2174), .B0(N2176));
NOR2XL inst_cellmath__24_0_I1171 (.Y(N2203), .A(N2177), .B(N2175));
OAI21XL inst_cellmath__24_0_I1172 (.Y(N2204), .A0(N2181), .A1(N2178), .B0(N2180));
NOR2XL inst_cellmath__24_0_I1173 (.Y(N2205), .A(N2181), .B(N2179));
OAI21XL inst_cellmath__24_0_I1174 (.Y(N2206), .A0(N2185), .A1(N2182), .B0(N2184));
NOR2XL inst_cellmath__24_0_I1175 (.Y(N2207), .A(N2185), .B(N2183));
OAI21XL inst_cellmath__24_0_I1176 (.Y(N2208), .A0(N2189), .A1(N2186), .B0(N2188));
NOR2XL inst_cellmath__24_0_I1177 (.Y(N2209), .A(N2189), .B(N2187));
OAI21XL inst_cellmath__24_0_I1178 (.Y(N2210), .A0(N2193), .A1(N2190), .B0(N2192));
NOR2XL inst_cellmath__24_0_I1179 (.Y(N2211), .A(N2193), .B(N2191));
AOI21XL inst_cellmath__24_0_I1182 (.Y(N2214), .A0(N2203), .A1(N2200), .B0(N2202));
AOI21XL inst_cellmath__24_0_I1184 (.Y(N2216), .A0(N2207), .A1(N2204), .B0(N2206));
NAND2XL inst_cellmath__24_0_I1185 (.Y(N2217), .A(N2207), .B(N2205));
AOI21XL inst_cellmath__24_0_I1186 (.Y(N2218), .A0(N2211), .A1(N2208), .B0(N2210));
OAI21XL inst_cellmath__24_0_I1188 (.Y(N2220), .A0(N2217), .A1(N2214), .B0(N2216));
INVXL inst_cellmath__24_0_I1190 (.Y(N2222), .A(N2205));
INVXL inst_cellmath__24_0_I1191 (.Y(N2223), .A(N2204));
OAI21XL inst_cellmath__24_0_I1192 (.Y(N2224), .A0(N2222), .A1(N2214), .B0(N2223));
INVXL inst_cellmath__24_0_I2477 (.Y(N7128), .A(N2220));
AOI21XL inst_cellmath__24_0_I1196 (.Y(N2228), .A0(N2209), .A1(N2220), .B0(N2208));
INVXL inst_cellmath__24_0_I1199 (.Y(N2231), .A(N2218));
AOI31X1 inst_cellmath__24_0_I2524 (.Y(N2232), .A0(N2211), .A1(N2209), .A2(N2220), .B0(N2231));
INVXL inst_cellmath__24_0_I1202 (.Y(N2234), .A(N2175));
INVXL inst_cellmath__24_0_I1203 (.Y(N2235), .A(N2174));
AOI21XL inst_cellmath__24_0_I1204 (.Y(N2236), .A0(N2234), .A1(N2200), .B0(N2235));
INVXL inst_cellmath__24_0_I2480 (.Y(N7131), .A(N2214));
OAI21XL inst_cellmath__24_0_I1208 (.Y(N2240), .A0(N2179), .A1(N2214), .B0(N2178));
INVXL inst_cellmath__24_0_I2481 (.Y(N7132), .A(N2224));
INVXL inst_cellmath__24_0_I1212 (.Y(N2244), .A(N2183));
INVXL inst_cellmath__24_0_I1213 (.Y(N2245), .A(N2182));
AOI21XL inst_cellmath__24_0_I1214 (.Y(N2246), .A0(N2244), .A1(N2224), .B0(N2245));
INVXL inst_cellmath__24_0_I2482 (.Y(N7133), .A(N7128));
OAI21XL inst_cellmath__24_0_I1218 (.Y(N2250), .A0(N2187), .A1(N7128), .B0(N2186));
INVXL inst_cellmath__24_0_I2483 (.Y(N7134), .A(N2228));
OAI21XL inst_cellmath__24_0_I1222 (.Y(N2254), .A0(N2191), .A1(N2228), .B0(N2190));
INVXL inst_cellmath__24_0_I2484 (.Y(N7135), .A(N2232));
OAI21XL inst_cellmath__24_0_I1226 (.Y(N2258), .A0(N2195), .A1(N2232), .B0(N2194));
OA21X1 inst_cellmath__24_0_I2254 (.Y(N2261), .A0(N2197), .A1(N2194), .B0(N2196));
OAI31X1 inst_cellmath__24_0_I2525 (.Y(N2262), .A0(N2197), .A1(N2195), .A2(N2232), .B0(N2261));
INVXL inst_cellmath__24_0_I1232 (.Y(N2264), .A(N2115));
INVXL inst_cellmath__24_0_I1233 (.Y(N2265), .A(N2114));
OAI21XL inst_cellmath__24_0_I1234 (.Y(N2266), .A0(N2264), .A1(N2170), .B0(N2265));
AOI21XL inst_cellmath__24_0_I1238 (.Y(N2270), .A0(N2119), .A1(N2200), .B0(N2118));
INVXL inst_cellmath__24_0_I1242 (.Y(N2274), .A(N2123));
INVXL inst_cellmath__24_0_I1243 (.Y(N2275), .A(N2122));
OAI21XL inst_cellmath__24_0_I1244 (.Y(N2276), .A0(N2274), .A1(N2236), .B0(N2275));
AOI21XL inst_cellmath__24_0_I1248 (.Y(N2280), .A0(N2127), .A1(N7131), .B0(N2126));
AOI21XL inst_cellmath__24_0_I1252 (.Y(N2284), .A0(N2131), .A1(N2240), .B0(N2130));
INVXL inst_cellmath__24_0_I1256 (.Y(N2288), .A(N2135));
INVXL inst_cellmath__24_0_I1257 (.Y(N2289), .A(N2134));
OAI21XL inst_cellmath__24_0_I1258 (.Y(N2290), .A0(N2288), .A1(N7132), .B0(N2289));
INVXL inst_cellmath__24_0_I1262 (.Y(N2294), .A(N2139));
INVXL inst_cellmath__24_0_I1263 (.Y(N2295), .A(N2138));
OAI21XL inst_cellmath__24_0_I1264 (.Y(N2296), .A0(N2294), .A1(N2246), .B0(N2295));
AOI21XL inst_cellmath__24_0_I1268 (.Y(N2300), .A0(N2143), .A1(N7133), .B0(N2142));
AOI21XL inst_cellmath__24_0_I1272 (.Y(N2304), .A0(N2147), .A1(N2250), .B0(N2146));
AOI21XL inst_cellmath__24_0_I1276 (.Y(N2308), .A0(N2151), .A1(N7134), .B0(N2150));
AOI21XL inst_cellmath__24_0_I1280 (.Y(N2312), .A0(N2155), .A1(N2254), .B0(N2154));
AOI21XL inst_cellmath__24_0_I1284 (.Y(N2316), .A0(N2159), .A1(N7135), .B0(N2158));
AOI21XL inst_cellmath__24_0_I1288 (.Y(N2320), .A0(N2163), .A1(N2258), .B0(N2162));
AOI21XL inst_cellmath__24_0_I1292 (.Y(N2324), .A0(N2167), .A1(N2262), .B0(N2166));
XNOR2X1 inst_cellmath__24_0_I1302 (.Y(inst_cellmath__24_0_out0[19]), .A(N2110), .B(N2113));
XOR2XL inst_cellmath__24_0_I1303 (.Y(inst_cellmath__24_0_out0[20]), .A(N2170), .B(N2115));
XNOR2X1 inst_cellmath__24_0_I1304 (.Y(inst_cellmath__24_0_out0[21]), .A(N2266), .B(N2117));
XNOR2X1 inst_cellmath__24_0_I1305 (.Y(inst_cellmath__24_0_out0[22]), .A(N2200), .B(N2119));
XOR2XL inst_cellmath__24_0_I1306 (.Y(inst_cellmath__24_0_out0[23]), .A(N2270), .B(N2121));
XOR2XL inst_cellmath__24_0_I2526 (.Y(inst_cellmath__24_0_out0[24]), .A(N2236), .B(N2123));
XNOR2X1 inst_cellmath__24_0_I1308 (.Y(inst_cellmath__24_0_out0[25]), .A(N2276), .B(N2125));
XNOR2X1 inst_cellmath__24_0_I1309 (.Y(inst_cellmath__24_0_out0[26]), .A(N7131), .B(N2127));
XOR2XL inst_cellmath__24_0_I1310 (.Y(inst_cellmath__24_0_out0[27]), .A(N2280), .B(N2129));
XNOR2X1 inst_cellmath__24_0_I1311 (.Y(inst_cellmath__24_0_out0[28]), .A(N2240), .B(N2131));
XOR2XL inst_cellmath__24_0_I1312 (.Y(inst_cellmath__24_0_out0[29]), .A(N2284), .B(N2133));
XOR2XL inst_cellmath__24_0_I2527 (.Y(inst_cellmath__24_0_out0[30]), .A(N7132), .B(N2135));
XNOR2X1 inst_cellmath__24_0_I1314 (.Y(inst_cellmath__24_0_out0[31]), .A(N2290), .B(N2137));
XOR2XL inst_cellmath__24_0_I2528 (.Y(inst_cellmath__24_0_out0[32]), .A(N2246), .B(N2139));
XNOR2X1 inst_cellmath__24_0_I1316 (.Y(inst_cellmath__24_0_out0[33]), .A(N2296), .B(N2141));
XNOR2X1 inst_cellmath__24_0_I1317 (.Y(inst_cellmath__24_0_out0[34]), .A(N7133), .B(N2143));
XOR2XL inst_cellmath__24_0_I1318 (.Y(inst_cellmath__24_0_out0[35]), .A(N2300), .B(N2145));
XNOR2X1 inst_cellmath__24_0_I1319 (.Y(inst_cellmath__24_0_out0[36]), .A(N2250), .B(N2147));
XOR2XL inst_cellmath__24_0_I1320 (.Y(inst_cellmath__24_0_out0[37]), .A(N2304), .B(N2149));
XNOR2X1 inst_cellmath__24_0_I1321 (.Y(inst_cellmath__24_0_out0[38]), .A(N7134), .B(N2151));
XOR2XL inst_cellmath__24_0_I1322 (.Y(inst_cellmath__24_0_out0[39]), .A(N2308), .B(N2153));
XNOR2X1 inst_cellmath__24_0_I1323 (.Y(inst_cellmath__24_0_out0[40]), .A(N2254), .B(N2155));
XOR2XL inst_cellmath__24_0_I1324 (.Y(inst_cellmath__24_0_out0[41]), .A(N2312), .B(N2157));
XNOR2X1 inst_cellmath__24_0_I1325 (.Y(inst_cellmath__24_0_out0[42]), .A(N7135), .B(N2159));
XOR2XL inst_cellmath__24_0_I1326 (.Y(inst_cellmath__24_0_out0[43]), .A(N2316), .B(N2161));
XNOR2X1 inst_cellmath__24_0_I1327 (.Y(inst_cellmath__24_0_out0[44]), .A(N2258), .B(N2163));
XOR2XL inst_cellmath__24_0_I1328 (.Y(inst_cellmath__24_0_out0[45]), .A(N2320), .B(N2165));
XNOR2X1 inst_cellmath__24_0_I1329 (.Y(inst_cellmath__24_0_out0[46]), .A(N2262), .B(N2167));
XNOR2X1 inst_cellmath__24_0_I1330 (.Y(inst_cellmath__24_0_out0[47]), .A(N2324), .B(N2169));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__25_0_bdw2052368036_bdw (
	inst_cellmath__25_0_out0,
	inst_cellmath__25_0_in0
	); /* architecture "gate_level" */ 
output [47:0] inst_cellmath__25_0_out0;
input [47:0] inst_cellmath__25_0_in0;
wire N199;
BUFX2 inst_cellmath__25_0_I51 (.Y(N199), .A(inst_cellmath__25_0_in0[47]));
AND2XL inst_cellmath__25_0_I0 (.Y(inst_cellmath__25_0_out0[0]), .A(N199), .B(inst_cellmath__25_0_in0[0]));
MX2XL inst_cellmath__25_0_I1 (.Y(inst_cellmath__25_0_out0[1]), .A(inst_cellmath__25_0_in0[0]), .B(inst_cellmath__25_0_in0[1]), .S0(N199));
MX2XL inst_cellmath__25_0_I2 (.Y(inst_cellmath__25_0_out0[2]), .A(inst_cellmath__25_0_in0[1]), .B(inst_cellmath__25_0_in0[2]), .S0(N199));
MX2XL inst_cellmath__25_0_I3 (.Y(inst_cellmath__25_0_out0[3]), .A(inst_cellmath__25_0_in0[2]), .B(inst_cellmath__25_0_in0[3]), .S0(N199));
MX2XL inst_cellmath__25_0_I4 (.Y(inst_cellmath__25_0_out0[4]), .A(inst_cellmath__25_0_in0[3]), .B(inst_cellmath__25_0_in0[4]), .S0(N199));
MX2XL inst_cellmath__25_0_I5 (.Y(inst_cellmath__25_0_out0[5]), .A(inst_cellmath__25_0_in0[4]), .B(inst_cellmath__25_0_in0[5]), .S0(N199));
MX2XL inst_cellmath__25_0_I6 (.Y(inst_cellmath__25_0_out0[6]), .A(inst_cellmath__25_0_in0[5]), .B(inst_cellmath__25_0_in0[6]), .S0(N199));
MX2XL inst_cellmath__25_0_I7 (.Y(inst_cellmath__25_0_out0[7]), .A(inst_cellmath__25_0_in0[6]), .B(inst_cellmath__25_0_in0[7]), .S0(N199));
MX2XL inst_cellmath__25_0_I8 (.Y(inst_cellmath__25_0_out0[8]), .A(inst_cellmath__25_0_in0[7]), .B(inst_cellmath__25_0_in0[8]), .S0(N199));
MX2XL inst_cellmath__25_0_I9 (.Y(inst_cellmath__25_0_out0[9]), .A(inst_cellmath__25_0_in0[8]), .B(inst_cellmath__25_0_in0[9]), .S0(N199));
MX2XL inst_cellmath__25_0_I10 (.Y(inst_cellmath__25_0_out0[10]), .A(inst_cellmath__25_0_in0[9]), .B(inst_cellmath__25_0_in0[10]), .S0(N199));
MX2XL inst_cellmath__25_0_I11 (.Y(inst_cellmath__25_0_out0[11]), .A(inst_cellmath__25_0_in0[10]), .B(inst_cellmath__25_0_in0[11]), .S0(N199));
MX2XL inst_cellmath__25_0_I12 (.Y(inst_cellmath__25_0_out0[12]), .A(inst_cellmath__25_0_in0[11]), .B(inst_cellmath__25_0_in0[12]), .S0(N199));
MX2XL inst_cellmath__25_0_I13 (.Y(inst_cellmath__25_0_out0[13]), .A(inst_cellmath__25_0_in0[12]), .B(inst_cellmath__25_0_in0[13]), .S0(N199));
MX2XL inst_cellmath__25_0_I14 (.Y(inst_cellmath__25_0_out0[14]), .A(inst_cellmath__25_0_in0[13]), .B(inst_cellmath__25_0_in0[14]), .S0(N199));
MX2XL inst_cellmath__25_0_I15 (.Y(inst_cellmath__25_0_out0[15]), .A(inst_cellmath__25_0_in0[14]), .B(inst_cellmath__25_0_in0[15]), .S0(N199));
MX2XL inst_cellmath__25_0_I16 (.Y(inst_cellmath__25_0_out0[16]), .A(inst_cellmath__25_0_in0[15]), .B(inst_cellmath__25_0_in0[16]), .S0(N199));
MX2XL inst_cellmath__25_0_I17 (.Y(inst_cellmath__25_0_out0[17]), .A(inst_cellmath__25_0_in0[16]), .B(inst_cellmath__25_0_in0[17]), .S0(N199));
MX2XL inst_cellmath__25_0_I18 (.Y(inst_cellmath__25_0_out0[18]), .A(inst_cellmath__25_0_in0[17]), .B(inst_cellmath__25_0_in0[18]), .S0(N199));
MX2XL inst_cellmath__25_0_I19 (.Y(inst_cellmath__25_0_out0[19]), .A(inst_cellmath__25_0_in0[18]), .B(inst_cellmath__25_0_in0[19]), .S0(N199));
MX2XL inst_cellmath__25_0_I20 (.Y(inst_cellmath__25_0_out0[20]), .A(inst_cellmath__25_0_in0[19]), .B(inst_cellmath__25_0_in0[20]), .S0(N199));
MX2XL inst_cellmath__25_0_I21 (.Y(inst_cellmath__25_0_out0[21]), .A(inst_cellmath__25_0_in0[20]), .B(inst_cellmath__25_0_in0[21]), .S0(N199));
MX2XL inst_cellmath__25_0_I22 (.Y(inst_cellmath__25_0_out0[22]), .A(inst_cellmath__25_0_in0[21]), .B(inst_cellmath__25_0_in0[22]), .S0(N199));
MX2XL inst_cellmath__25_0_I23 (.Y(inst_cellmath__25_0_out0[23]), .A(inst_cellmath__25_0_in0[22]), .B(inst_cellmath__25_0_in0[23]), .S0(N199));
MX2XL inst_cellmath__25_0_I24 (.Y(inst_cellmath__25_0_out0[24]), .A(inst_cellmath__25_0_in0[23]), .B(inst_cellmath__25_0_in0[24]), .S0(N199));
MX2XL inst_cellmath__25_0_I25 (.Y(inst_cellmath__25_0_out0[25]), .A(inst_cellmath__25_0_in0[24]), .B(inst_cellmath__25_0_in0[25]), .S0(N199));
MX2XL inst_cellmath__25_0_I26 (.Y(inst_cellmath__25_0_out0[26]), .A(inst_cellmath__25_0_in0[25]), .B(inst_cellmath__25_0_in0[26]), .S0(N199));
MX2XL inst_cellmath__25_0_I27 (.Y(inst_cellmath__25_0_out0[27]), .A(inst_cellmath__25_0_in0[26]), .B(inst_cellmath__25_0_in0[27]), .S0(N199));
MX2XL inst_cellmath__25_0_I28 (.Y(inst_cellmath__25_0_out0[28]), .A(inst_cellmath__25_0_in0[27]), .B(inst_cellmath__25_0_in0[28]), .S0(N199));
MX2XL inst_cellmath__25_0_I29 (.Y(inst_cellmath__25_0_out0[29]), .A(inst_cellmath__25_0_in0[28]), .B(inst_cellmath__25_0_in0[29]), .S0(N199));
MX2XL inst_cellmath__25_0_I30 (.Y(inst_cellmath__25_0_out0[30]), .A(inst_cellmath__25_0_in0[29]), .B(inst_cellmath__25_0_in0[30]), .S0(N199));
MX2XL inst_cellmath__25_0_I31 (.Y(inst_cellmath__25_0_out0[31]), .A(inst_cellmath__25_0_in0[30]), .B(inst_cellmath__25_0_in0[31]), .S0(N199));
MX2XL inst_cellmath__25_0_I32 (.Y(inst_cellmath__25_0_out0[32]), .A(inst_cellmath__25_0_in0[31]), .B(inst_cellmath__25_0_in0[32]), .S0(N199));
MX2XL inst_cellmath__25_0_I33 (.Y(inst_cellmath__25_0_out0[33]), .A(inst_cellmath__25_0_in0[32]), .B(inst_cellmath__25_0_in0[33]), .S0(N199));
MX2XL inst_cellmath__25_0_I34 (.Y(inst_cellmath__25_0_out0[34]), .A(inst_cellmath__25_0_in0[33]), .B(inst_cellmath__25_0_in0[34]), .S0(N199));
MX2XL inst_cellmath__25_0_I35 (.Y(inst_cellmath__25_0_out0[35]), .A(inst_cellmath__25_0_in0[34]), .B(inst_cellmath__25_0_in0[35]), .S0(N199));
MX2XL inst_cellmath__25_0_I36 (.Y(inst_cellmath__25_0_out0[36]), .A(inst_cellmath__25_0_in0[35]), .B(inst_cellmath__25_0_in0[36]), .S0(N199));
MX2XL inst_cellmath__25_0_I37 (.Y(inst_cellmath__25_0_out0[37]), .A(inst_cellmath__25_0_in0[36]), .B(inst_cellmath__25_0_in0[37]), .S0(N199));
MX2XL inst_cellmath__25_0_I38 (.Y(inst_cellmath__25_0_out0[38]), .A(inst_cellmath__25_0_in0[37]), .B(inst_cellmath__25_0_in0[38]), .S0(N199));
MX2XL inst_cellmath__25_0_I39 (.Y(inst_cellmath__25_0_out0[39]), .A(inst_cellmath__25_0_in0[38]), .B(inst_cellmath__25_0_in0[39]), .S0(N199));
MX2XL inst_cellmath__25_0_I40 (.Y(inst_cellmath__25_0_out0[40]), .A(inst_cellmath__25_0_in0[39]), .B(inst_cellmath__25_0_in0[40]), .S0(N199));
MX2XL inst_cellmath__25_0_I41 (.Y(inst_cellmath__25_0_out0[41]), .A(inst_cellmath__25_0_in0[40]), .B(inst_cellmath__25_0_in0[41]), .S0(N199));
MX2XL inst_cellmath__25_0_I42 (.Y(inst_cellmath__25_0_out0[42]), .A(inst_cellmath__25_0_in0[41]), .B(inst_cellmath__25_0_in0[42]), .S0(N199));
MX2XL inst_cellmath__25_0_I43 (.Y(inst_cellmath__25_0_out0[43]), .A(inst_cellmath__25_0_in0[42]), .B(inst_cellmath__25_0_in0[43]), .S0(N199));
MX2XL inst_cellmath__25_0_I44 (.Y(inst_cellmath__25_0_out0[44]), .A(inst_cellmath__25_0_in0[43]), .B(inst_cellmath__25_0_in0[44]), .S0(N199));
MX2XL inst_cellmath__25_0_I45 (.Y(inst_cellmath__25_0_out0[45]), .A(inst_cellmath__25_0_in0[44]), .B(inst_cellmath__25_0_in0[45]), .S0(N199));
MX2XL inst_cellmath__25_0_I46 (.Y(inst_cellmath__25_0_out0[46]), .A(inst_cellmath__25_0_in0[45]), .B(inst_cellmath__25_0_in0[46]), .S0(N199));
OR2XL inst_cellmath__25_0_I47 (.Y(inst_cellmath__25_0_out0[47]), .A(N199), .B(inst_cellmath__25_0_in0[46]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__45_0_bdw2052368036_bdw (
	inst_cellmath__45_0_out0,
	inst_cellmath__45_0_in0
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__45_0_out0;
input [47:24] inst_cellmath__45_0_in0;
wire N146,N154,N160,N164,N172,N181,N184 
	,N187,N190,N196,N200,N208,N212,N216,N224 
	,N238,N240,N263,N272,N278,N284,N288,N296 
	,N300,N312,N328,N381,N384,N387,N390,N393 
	,N396,N399,N402,N733,N743,N749,N750,N752 
	,N753,N755,N763;
INVXL inst_cellmath__45_0_I37 (.Y(inst_cellmath__45_0_out0[0]), .A(inst_cellmath__45_0_in0[24]));
NAND2XL inst_cellmath__45_0_I42 (.Y(N146), .A(inst_cellmath__45_0_in0[26]), .B(inst_cellmath__45_0_in0[25]));
NOR2XL inst_cellmath__45_0_I49 (.Y(N154), .A(N146), .B(inst_cellmath__45_0_out0[0]));
NAND2XL inst_cellmath__45_0_I54 (.Y(N160), .A(inst_cellmath__45_0_in0[28]), .B(inst_cellmath__45_0_in0[27]));
NAND2XL inst_cellmath__45_0_I58 (.Y(N164), .A(inst_cellmath__45_0_in0[30]), .B(inst_cellmath__45_0_in0[29]));
NOR2XL inst_cellmath__45_0_I66 (.Y(N172), .A(N164), .B(N160));
NAND2XL inst_cellmath__45_0_I75 (.Y(N181), .A(inst_cellmath__45_0_in0[27]), .B(N154));
NAND2BXL inst_cellmath__45_0_I565 (.Y(N184), .AN(N160), .B(N154));
NAND3BXL inst_cellmath__45_0_I566 (.Y(N187), .AN(N160), .B(inst_cellmath__45_0_in0[29]), .C(N154));
NAND2XL inst_cellmath__45_0_I81 (.Y(N190), .A(N172), .B(N154));
NAND2XL inst_cellmath__45_0_I86 (.Y(N196), .A(inst_cellmath__45_0_in0[32]), .B(inst_cellmath__45_0_in0[31]));
NAND2XL inst_cellmath__45_0_I90 (.Y(N200), .A(inst_cellmath__45_0_in0[34]), .B(inst_cellmath__45_0_in0[33]));
NOR2XL inst_cellmath__45_0_I98 (.Y(N208), .A(N200), .B(N196));
NAND2XL inst_cellmath__45_0_I102 (.Y(N212), .A(inst_cellmath__45_0_in0[36]), .B(inst_cellmath__45_0_in0[35]));
NAND2XL inst_cellmath__45_0_I106 (.Y(N216), .A(inst_cellmath__45_0_in0[38]), .B(inst_cellmath__45_0_in0[37]));
NOR2XL inst_cellmath__45_0_I114 (.Y(N224), .A(N216), .B(N212));
NAND3BXL inst_cellmath__45_0_I575 (.Y(N238), .AN(N212), .B(inst_cellmath__45_0_in0[37]), .C(N208));
NAND2XL inst_cellmath__45_0_I130 (.Y(N240), .A(N224), .B(N208));
NOR3BXL inst_cellmath__45_0_I577 (.Y(N263), .AN(inst_cellmath__45_0_in0[33]), .B(N196), .C(N190));
NOR3BXL inst_cellmath__45_0_I579 (.Y(N272), .AN(N208), .B(N212), .C(N190));
NOR2XL inst_cellmath__45_0_I161 (.Y(N278), .A(N240), .B(N190));
NAND2XL inst_cellmath__45_0_I166 (.Y(N284), .A(inst_cellmath__45_0_in0[40]), .B(inst_cellmath__45_0_in0[39]));
NAND2XL inst_cellmath__45_0_I170 (.Y(N288), .A(inst_cellmath__45_0_in0[42]), .B(inst_cellmath__45_0_in0[41]));
NOR2XL inst_cellmath__45_0_I178 (.Y(N296), .A(N288), .B(N284));
NAND2XL inst_cellmath__45_0_I182 (.Y(N300), .A(inst_cellmath__45_0_in0[44]), .B(inst_cellmath__45_0_in0[43]));
NAND2XL hyperpropagate_3_1_A_I627 (.Y(N763), .A(inst_cellmath__45_0_in0[46]), .B(inst_cellmath__45_0_in0[45]));
NOR2XL hyperpropagate_3_1_A_I628 (.Y(N312), .A(N300), .B(N763));
NAND2XL inst_cellmath__45_0_I210 (.Y(N328), .A(N312), .B(N296));
INVXL inst_cellmath__45_0_I531 (.Y(N733), .A(inst_cellmath__45_0_in0[47]));
NAND2BXL inst_cellmath__45_0_I593 (.Y(N743), .AN(inst_cellmath__45_0_out0[0]), .B(inst_cellmath__45_0_in0[25]));
NAND2BXL inst_cellmath__45_0_I594 (.Y(N749), .AN(N190), .B(inst_cellmath__45_0_in0[31]));
OR2XL inst_cellmath__45_0_I595 (.Y(N750), .A(N196), .B(N190));
NAND2BXL inst_cellmath__45_0_I596 (.Y(N752), .AN(N190), .B(N208));
NAND3BXL inst_cellmath__45_0_I616 (.Y(N753), .AN(N190), .B(inst_cellmath__45_0_in0[35]), .C(N208));
OR2XL inst_cellmath__45_0_I598 (.Y(N755), .A(N238), .B(N190));
NAND2XL inst_cellmath__45_0_I263 (.Y(N381), .A(inst_cellmath__45_0_in0[39]), .B(N278));
NAND2BXL inst_cellmath__45_0_I599 (.Y(N384), .AN(N284), .B(N278));
NAND3BXL inst_cellmath__45_0_I600 (.Y(N387), .AN(N284), .B(inst_cellmath__45_0_in0[41]), .C(N278));
NAND2XL inst_cellmath__45_0_I269 (.Y(N390), .A(N296), .B(N278));
NAND3XL inst_cellmath__45_0_I601 (.Y(N393), .A(inst_cellmath__45_0_in0[43]), .B(N296), .C(N278));
NAND3BXL inst_cellmath__45_0_I602 (.Y(N396), .AN(N300), .B(N296), .C(N278));
NAND4BXL inst_cellmath__45_0_I603 (.Y(N399), .AN(N300), .B(inst_cellmath__45_0_in0[45]), .C(N278), .D(N296));
NAND2BXL inst_cellmath__45_0_I604 (.Y(N402), .AN(N328), .B(N278));
NOR3BXL inst_cellmath__45_0_I767 (.Y(inst_cellmath__45_0_out0[24]), .AN(N278), .B(N733), .C(N328));
XNOR2X1 inst_cellmath__45_0_I380 (.Y(inst_cellmath__45_0_out0[1]), .A(inst_cellmath__45_0_out0[0]), .B(inst_cellmath__45_0_in0[25]));
XNOR2X1 inst_cellmath__45_0_I381 (.Y(inst_cellmath__45_0_out0[2]), .A(N743), .B(inst_cellmath__45_0_in0[26]));
XOR2XL inst_cellmath__45_0_I606 (.Y(inst_cellmath__45_0_out0[3]), .A(N154), .B(inst_cellmath__45_0_in0[27]));
XNOR2X1 inst_cellmath__45_0_I383 (.Y(inst_cellmath__45_0_out0[4]), .A(N181), .B(inst_cellmath__45_0_in0[28]));
XNOR2X1 inst_cellmath__45_0_I384 (.Y(inst_cellmath__45_0_out0[5]), .A(N184), .B(inst_cellmath__45_0_in0[29]));
XNOR2X1 inst_cellmath__45_0_I385 (.Y(inst_cellmath__45_0_out0[6]), .A(N187), .B(inst_cellmath__45_0_in0[30]));
XNOR2X1 inst_cellmath__45_0_I386 (.Y(inst_cellmath__45_0_out0[7]), .A(N190), .B(inst_cellmath__45_0_in0[31]));
XNOR2X1 inst_cellmath__45_0_I387 (.Y(inst_cellmath__45_0_out0[8]), .A(N749), .B(inst_cellmath__45_0_in0[32]));
XNOR2X1 inst_cellmath__45_0_I388 (.Y(inst_cellmath__45_0_out0[9]), .A(N750), .B(inst_cellmath__45_0_in0[33]));
XOR2XL inst_cellmath__45_0_I607 (.Y(inst_cellmath__45_0_out0[10]), .A(N263), .B(inst_cellmath__45_0_in0[34]));
XNOR2X1 inst_cellmath__45_0_I390 (.Y(inst_cellmath__45_0_out0[11]), .A(N752), .B(inst_cellmath__45_0_in0[35]));
XNOR2X1 inst_cellmath__45_0_I391 (.Y(inst_cellmath__45_0_out0[12]), .A(N753), .B(inst_cellmath__45_0_in0[36]));
XOR2XL inst_cellmath__45_0_I608 (.Y(inst_cellmath__45_0_out0[13]), .A(N272), .B(inst_cellmath__45_0_in0[37]));
XNOR2X1 inst_cellmath__45_0_I393 (.Y(inst_cellmath__45_0_out0[14]), .A(N755), .B(inst_cellmath__45_0_in0[38]));
XOR2XL inst_cellmath__45_0_I609 (.Y(inst_cellmath__45_0_out0[15]), .A(N278), .B(inst_cellmath__45_0_in0[39]));
XNOR2X1 inst_cellmath__45_0_I395 (.Y(inst_cellmath__45_0_out0[16]), .A(N381), .B(inst_cellmath__45_0_in0[40]));
XNOR2X1 inst_cellmath__45_0_I396 (.Y(inst_cellmath__45_0_out0[17]), .A(N384), .B(inst_cellmath__45_0_in0[41]));
XNOR2X1 inst_cellmath__45_0_I397 (.Y(inst_cellmath__45_0_out0[18]), .A(N387), .B(inst_cellmath__45_0_in0[42]));
XNOR2X1 inst_cellmath__45_0_I398 (.Y(inst_cellmath__45_0_out0[19]), .A(N390), .B(inst_cellmath__45_0_in0[43]));
XNOR2X1 inst_cellmath__45_0_I399 (.Y(inst_cellmath__45_0_out0[20]), .A(N393), .B(inst_cellmath__45_0_in0[44]));
XNOR2X1 inst_cellmath__45_0_I400 (.Y(inst_cellmath__45_0_out0[21]), .A(N396), .B(inst_cellmath__45_0_in0[45]));
XNOR2X1 inst_cellmath__45_0_I401 (.Y(inst_cellmath__45_0_out0[22]), .A(N399), .B(inst_cellmath__45_0_in0[46]));
XOR2XL inst_cellmath__45_0_I610 (.Y(inst_cellmath__45_0_out0[23]), .A(N733), .B(N402));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__5_1_bdw2052368036_bdw (
	inst_cellmath__5_1_out0,
	inst_cellmath__5_1_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__5_1_out0;
input [2:0] inst_cellmath__5_1_in0;
NOR3BXL inst_cellmath__5_1_I17 (.Y(inst_cellmath__5_1_out0), .AN(inst_cellmath__5_1_in0[0]), .B(inst_cellmath__5_1_in0[2]), .C(inst_cellmath__5_1_in0[1]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__31__bdw2052368036_bdw (
	inst_cellmath__44__31__out0,
	inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__31__out0;
input  inst_cellmath__44__31__in0,
	inst_cellmath__44__31__in1;
wire N13;
INVXL inst_cellmath__44__31__I3 (.Y(N13), .A(inst_cellmath__44__31__in1));
AND2XL inst_cellmath__44__31__I1 (.Y(inst_cellmath__44__31__out0[0]), .A(inst_cellmath__44__31__in0), .B(N13));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__6_0_bdw2052368036_bdw (
	inst_cellmath__6_0_out0,
	inst_cellmath__6_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__6_0_out0;
input [2:0] inst_cellmath__6_0_in0;
NOR3BXL inst_cellmath__6_0_I23 (.Y(inst_cellmath__6_0_out0), .AN(inst_cellmath__6_0_in0[1]), .B(inst_cellmath__6_0_in0[2]), .C(inst_cellmath__6_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__30__bdw2052368036_bdw (
	inst_cellmath__44__30__out0,
	inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__30__out0;
input  inst_cellmath__44__30__in0,
	inst_cellmath__44__30__in1;
AND2XL inst_cellmath__44__30__I0 (.Y(inst_cellmath__44__30__out0[0]), .A(inst_cellmath__44__30__in0), .B(inst_cellmath__44__30__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__8_0_bdw2052368036_bdw (
	inst_cellmath__8_0_out0,
	inst_cellmath__8_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__8_0_out0;
input [2:0] inst_cellmath__8_0_in0;
NOR3BXL inst_cellmath__8_0_I34 (.Y(inst_cellmath__8_0_out0), .AN(inst_cellmath__8_0_in0[2]), .B(inst_cellmath__8_0_in0[1]), .C(inst_cellmath__8_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__4_0_bdw2052368036_bdw (
	inst_cellmath__4_0_out0,
	inst_cellmath__4_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__4_0_out0;
input [2:0] inst_cellmath__4_0_in0;
NOR3XL inst_cellmath__4_0_I39 (.Y(inst_cellmath__4_0_out0), .A(inst_cellmath__4_0_in0[1]), .B(inst_cellmath__4_0_in0[2]), .C(inst_cellmath__4_0_in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__34_0_bdw2052368036_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__34_0_out0;
input [22:0] inst_cellmath__34_0_in0;
wire N29,N30,N31,N32,N33,N34,N35 
	,N36,N37,N38,N39,N40,N42,N43,N45 
	,N48,N49,N70;
NOR2XL inst_cellmath__34_0_I3 (.Y(N29), .A(inst_cellmath__34_0_in0[19]), .B(inst_cellmath__34_0_in0[17]));
NOR2XL inst_cellmath__34_0_I4 (.Y(N30), .A(inst_cellmath__34_0_in0[15]), .B(inst_cellmath__34_0_in0[13]));
NOR2XL inst_cellmath__34_0_I5 (.Y(N31), .A(inst_cellmath__34_0_in0[11]), .B(inst_cellmath__34_0_in0[9]));
NOR2XL inst_cellmath__34_0_I6 (.Y(N32), .A(inst_cellmath__34_0_in0[7]), .B(inst_cellmath__34_0_in0[5]));
NOR2XL inst_cellmath__34_0_I7 (.Y(N33), .A(inst_cellmath__34_0_in0[3]), .B(inst_cellmath__34_0_in0[22]));
NOR2XL inst_cellmath__34_0_I8 (.Y(N34), .A(inst_cellmath__34_0_in0[20]), .B(inst_cellmath__34_0_in0[18]));
NOR2XL inst_cellmath__34_0_I9 (.Y(N35), .A(inst_cellmath__34_0_in0[16]), .B(inst_cellmath__34_0_in0[14]));
NOR2XL inst_cellmath__34_0_I10 (.Y(N36), .A(inst_cellmath__34_0_in0[12]), .B(inst_cellmath__34_0_in0[10]));
NOR2XL inst_cellmath__34_0_I11 (.Y(N37), .A(inst_cellmath__34_0_in0[8]), .B(inst_cellmath__34_0_in0[6]));
NOR2XL inst_cellmath__34_0_I12 (.Y(N38), .A(inst_cellmath__34_0_in0[4]), .B(inst_cellmath__34_0_in0[2]));
NAND2XL inst_cellmath__34_0_I13 (.Y(N39), .A(N29), .B(N30));
NAND2XL inst_cellmath__34_0_I14 (.Y(N40), .A(N31), .B(N32));
NAND2XL inst_cellmath__34_0_I16 (.Y(N42), .A(N35), .B(N36));
NAND2XL inst_cellmath__34_0_I17 (.Y(N43), .A(N37), .B(N38));
NOR4X1 inst_cellmath__34_0_I27 (.Y(N45), .A(inst_cellmath__34_0_in0[0]), .B(inst_cellmath__34_0_in0[1]), .C(inst_cellmath__34_0_in0[21]), .D(N39));
NOR2XL inst_cellmath__34_0_I21 (.Y(N49), .A(N42), .B(N43));
NAND3XL hyperpropagate_4_1_A_I30 (.Y(N70), .A(N33), .B(N34), .C(N45));
NOR2XL hyperpropagate_4_1_A_I31 (.Y(N48), .A(N40), .B(N70));
NAND2XL inst_cellmath__34_0_I24 (.Y(inst_cellmath__34_0_out0), .A(N49), .B(N48));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__29__bdw2052368036_bdw (
	inst_cellmath__44__29__out0,
	inst_cellmath__44__29__in0,
	inst_cellmath__44__29__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__29__out0;
input  inst_cellmath__44__29__in0;
input [24:24] inst_cellmath__44__29__in1;
OR2XL inst_cellmath__44__29__I0 (.Y(inst_cellmath__44__29__out0[0]), .A(inst_cellmath__44__29__in1[24]), .B(inst_cellmath__44__29__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__28__bdw2052368036_bdw (
	inst_cellmath__44__28__out0,
	inst_cellmath__44__28__in0,
	inst_cellmath__44__28__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__28__out0;
input [0:0] inst_cellmath__44__28__in0;
input  inst_cellmath__44__28__in1;
AND2XL inst_cellmath__44__28__I0 (.Y(inst_cellmath__44__28__out0[0]), .A(inst_cellmath__44__28__in1), .B(inst_cellmath__44__28__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__27__bdw2052368036_bdw (
	inst_cellmath__44__27__out0,
	inst_cellmath__44__27__in0,
	inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__27__out0;
input  inst_cellmath__44__27__in0;
input [0:0] inst_cellmath__44__27__in1,
	inst_cellmath__44__27__in2,
	inst_cellmath__44__27__in3;
OR4X1 inst_cellmath__44__27__I7 (.Y(inst_cellmath__44__27__out0[0]), .A(inst_cellmath__44__27__in0), .B(inst_cellmath__44__27__in2[0]), .C(inst_cellmath__44__27__in1[0]), .D(inst_cellmath__44__27__in3[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__26__bdw2052368036_bdw (
	inst_cellmath__44__26__out0,
	inst_cellmath__44__26__in0,
	inst_cellmath__44__26__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__26__out0;
input [0:0] inst_cellmath__44__26__in0;
input [23:23] inst_cellmath__44__26__in1;
AND2XL inst_cellmath__44__26__I0 (.Y(inst_cellmath__44__26__out0[0]), .A(inst_cellmath__44__26__in1[23]), .B(inst_cellmath__44__26__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__33__bdw2052368036_bdw (
	inst_cellmath__44__33__out0,
	inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__33__out0;
input [0:0] inst_cellmath__44__33__in0,
	inst_cellmath__44__33__in1;
OR2XL inst_cellmath__44__33__I0 (.Y(inst_cellmath__44__33__out0[0]), .A(inst_cellmath__44__33__in1[0]), .B(inst_cellmath__44__33__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44__32__bdw2052368036_bdw (
	inst_cellmath__44__32__out0,
	inst_cellmath__44__32__in0,
	inst_cellmath__44__32__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__44__32__out0;
input [0:0] inst_cellmath__44__32__in0;
input  inst_cellmath__44__32__in1;
AND2XL inst_cellmath__44__32__I0 (.Y(inst_cellmath__44__32__out0[0]), .A(inst_cellmath__44__32__in0[0]), .B(inst_cellmath__44__32__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__44_0_bdw2052368036_bdw (
	inst_cellmath__44_0_out0,
	inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__44_0_out0;
input [0:0] inst_cellmath__44_0_in0,
	inst_cellmath__44_0_in1;
OR2XL inst_cellmath__44_0_I0 (.Y(inst_cellmath__44_0_out0), .A(inst_cellmath__44_0_in0[0]), .B(inst_cellmath__44_0_in1[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__46_0_bdw2052368036_bdw (
	inst_cellmath__46_0_out0,
	inst_cellmath__46_0_in0,
	inst_cellmath__46_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__46_0_out0;
input [24:24] inst_cellmath__46_0_in0;
input  inst_cellmath__46_0_in1;
AND2XL inst_cellmath__46_0_I0 (.Y(inst_cellmath__46_0_out0), .A(inst_cellmath__46_0_in0[24]), .B(inst_cellmath__46_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__38_0_bdw2052368036_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0;
input [47:47] inst_cellmath__38_0_in1;
OR2XL inst_cellmath__38_0_I0 (.Y(inst_cellmath__38_0_out0), .A(inst_cellmath__38_0_in1[47]), .B(inst_cellmath__38_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__30_0_bdw2052368036_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__30_0_out0;
input [7:0] inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
wire N106,N111,N115,N117,N119,N121,N123 
	,N125,N127;
INVXL inst_cellmath__30_0_I40 (.Y(N106), .A(inst_cellmath__30_0_in1[7]));
XNOR2X1 hap1_A_I51 (.Y(inst_cellmath__30_0_out0[0]), .A(inst_cellmath__30_0_in0[0]), .B(inst_cellmath__30_0_in1[0]));
OR2XL hap1_A_I52 (.Y(N111), .A(inst_cellmath__30_0_in0[0]), .B(inst_cellmath__30_0_in1[0]));
ADDFX1 inst_cellmath__30_0_I42 (.CO(N115), .S(inst_cellmath__30_0_out0[1]), .A(inst_cellmath__30_0_in0[1]), .B(inst_cellmath__30_0_in1[1]), .CI(N111));
ADDFX1 inst_cellmath__30_0_I43 (.CO(N117), .S(inst_cellmath__30_0_out0[2]), .A(inst_cellmath__30_0_in0[2]), .B(inst_cellmath__30_0_in1[2]), .CI(N115));
ADDFX1 inst_cellmath__30_0_I44 (.CO(N119), .S(inst_cellmath__30_0_out0[3]), .A(inst_cellmath__30_0_in0[3]), .B(inst_cellmath__30_0_in1[3]), .CI(N117));
ADDFX1 inst_cellmath__30_0_I45 (.CO(N121), .S(inst_cellmath__30_0_out0[4]), .A(inst_cellmath__30_0_in0[4]), .B(inst_cellmath__30_0_in1[4]), .CI(N119));
ADDFX1 inst_cellmath__30_0_I46 (.CO(N123), .S(inst_cellmath__30_0_out0[5]), .A(inst_cellmath__30_0_in0[5]), .B(inst_cellmath__30_0_in1[5]), .CI(N121));
ADDFX1 inst_cellmath__30_0_I47 (.CO(N125), .S(inst_cellmath__30_0_out0[6]), .A(inst_cellmath__30_0_in0[6]), .B(inst_cellmath__30_0_in1[6]), .CI(N123));
ADDFX1 inst_cellmath__30_0_I48 (.CO(N127), .S(inst_cellmath__30_0_out0[7]), .A(N106), .B(inst_cellmath__30_0_in0[7]), .CI(N125));
XNOR2X1 hap1_A_I53 (.Y(inst_cellmath__30_0_out0[8]), .A(inst_cellmath__30_0_in1[7]), .B(N127));
NOR2XL hap1_A_I54 (.Y(inst_cellmath__30_0_out0[9]), .A(inst_cellmath__30_0_in1[7]), .B(N127));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__31_0_bdw2052368036_bdw (
	inst_cellmath__31_0_out0,
	inst_cellmath__31_0_in0
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__31_0_out0;
input [9:0] inst_cellmath__31_0_in0;
wire N77,N116,N119,N128,N131,N134,N137 
	,N140;
INVXL inst_cellmath__31_0_I99 (.Y(inst_cellmath__31_0_out0[0]), .A(inst_cellmath__31_0_in0[0]));
NOR2BX1 inst_cellmath__31_0_I102 (.Y(N77), .AN(inst_cellmath__31_0_in0[1]), .B(inst_cellmath__31_0_out0[0]));
AND2XL inst_cellmath__31_0_I38 (.Y(N116), .A(inst_cellmath__31_0_in0[2]), .B(N77));
XNOR2X1 inst_cellmath__31_0_I55 (.Y(inst_cellmath__31_0_out0[1]), .A(inst_cellmath__31_0_out0[0]), .B(inst_cellmath__31_0_in0[1]));
XOR2XL inst_cellmath__31_0_I103 (.Y(inst_cellmath__31_0_out0[2]), .A(N77), .B(inst_cellmath__31_0_in0[2]));
AND2XL inst_cellmath__31_0_I60 (.Y(N119), .A(inst_cellmath__31_0_in0[3]), .B(N116));
AND3XL inst_cellmath__31_0_I104 (.Y(N128), .A(inst_cellmath__31_0_in0[4]), .B(inst_cellmath__31_0_in0[5]), .C(N119));
AND3XL inst_cellmath__31_0_I105 (.Y(N131), .A(inst_cellmath__31_0_in0[6]), .B(inst_cellmath__31_0_in0[7]), .C(N128));
NAND2XL inst_cellmath__31_0_I72 (.Y(N134), .A(inst_cellmath__31_0_in0[4]), .B(N119));
NAND2XL inst_cellmath__31_0_I74 (.Y(N137), .A(inst_cellmath__31_0_in0[6]), .B(N128));
NAND2XL inst_cellmath__31_0_I76 (.Y(N140), .A(inst_cellmath__31_0_in0[8]), .B(N131));
XOR2XL inst_cellmath__31_0_I84 (.Y(inst_cellmath__31_0_out0[3]), .A(N116), .B(inst_cellmath__31_0_in0[3]));
XOR2XL inst_cellmath__31_0_I85 (.Y(inst_cellmath__31_0_out0[4]), .A(N119), .B(inst_cellmath__31_0_in0[4]));
XNOR2X1 inst_cellmath__31_0_I86 (.Y(inst_cellmath__31_0_out0[5]), .A(N134), .B(inst_cellmath__31_0_in0[5]));
XOR2XL inst_cellmath__31_0_I87 (.Y(inst_cellmath__31_0_out0[6]), .A(N128), .B(inst_cellmath__31_0_in0[6]));
XNOR2X1 inst_cellmath__31_0_I88 (.Y(inst_cellmath__31_0_out0[7]), .A(N137), .B(inst_cellmath__31_0_in0[7]));
XOR2XL inst_cellmath__31_0_I89 (.Y(inst_cellmath__31_0_out0[8]), .A(N131), .B(inst_cellmath__31_0_in0[8]));
XNOR2X1 inst_cellmath__31_0_I90 (.Y(inst_cellmath__31_0_out0[9]), .A(N140), .B(inst_cellmath__31_0_in0[9]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__48_0_bdw2052368036_bdw (
	inst_cellmath__48_0_out0,
	inst_cellmath__48_0_in0,
	inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2
	); /* architecture "gate_level" */ 
output [9:0] inst_cellmath__48_0_out0;
input  inst_cellmath__48_0_in0;
input [9:0] inst_cellmath__48_0_in1,
	inst_cellmath__48_0_in2;
MX2XL inst_cellmath__48_0_I20 (.Y(inst_cellmath__48_0_out0[0]), .A(inst_cellmath__48_0_in2[0]), .B(inst_cellmath__48_0_in1[0]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I21 (.Y(inst_cellmath__48_0_out0[1]), .A(inst_cellmath__48_0_in2[1]), .B(inst_cellmath__48_0_in1[1]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I22 (.Y(inst_cellmath__48_0_out0[2]), .A(inst_cellmath__48_0_in2[2]), .B(inst_cellmath__48_0_in1[2]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I23 (.Y(inst_cellmath__48_0_out0[3]), .A(inst_cellmath__48_0_in2[3]), .B(inst_cellmath__48_0_in1[3]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I24 (.Y(inst_cellmath__48_0_out0[4]), .A(inst_cellmath__48_0_in2[4]), .B(inst_cellmath__48_0_in1[4]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I25 (.Y(inst_cellmath__48_0_out0[5]), .A(inst_cellmath__48_0_in2[5]), .B(inst_cellmath__48_0_in1[5]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I26 (.Y(inst_cellmath__48_0_out0[6]), .A(inst_cellmath__48_0_in2[6]), .B(inst_cellmath__48_0_in1[6]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I27 (.Y(inst_cellmath__48_0_out0[7]), .A(inst_cellmath__48_0_in2[7]), .B(inst_cellmath__48_0_in1[7]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I28 (.Y(inst_cellmath__48_0_out0[8]), .A(inst_cellmath__48_0_in2[8]), .B(inst_cellmath__48_0_in1[8]), .S0(inst_cellmath__48_0_in0));
MX2XL inst_cellmath__48_0_I29 (.Y(inst_cellmath__48_0_out0[9]), .A(inst_cellmath__48_0_in2[9]), .B(inst_cellmath__48_0_in1[9]), .S0(inst_cellmath__48_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__49__bdw2052368036_bdw (
	inst_cellmath__51__49__out0,
	inst_cellmath__51__49__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__49__out0;
input [7:0] inst_cellmath__51__49__in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__51__49__I0 (.Y(N11), .A(inst_cellmath__51__49__in0[1]), .B(inst_cellmath__51__49__in0[6]));
NAND2XL inst_cellmath__51__49__I1 (.Y(N12), .A(inst_cellmath__51__49__in0[0]), .B(inst_cellmath__51__49__in0[5]));
NAND2XL inst_cellmath__51__49__I2 (.Y(N13), .A(inst_cellmath__51__49__in0[4]), .B(inst_cellmath__51__49__in0[2]));
NAND2XL inst_cellmath__51__49__I3 (.Y(N14), .A(inst_cellmath__51__49__in0[7]), .B(inst_cellmath__51__49__in0[3]));
NOR2XL inst_cellmath__51__49__I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__51__49__I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__51__49__I6 (.Y(inst_cellmath__51__49__out0[0]), .A(N15), .B(N16));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51__48__bdw2052368036_bdw (
	inst_cellmath__51__48__out0,
	inst_cellmath__51__48__in0,
	inst_cellmath__51__48__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__51__48__out0;
input [0:0] inst_cellmath__51__48__in0;
input [8:8] inst_cellmath__51__48__in1;
OR2XL inst_cellmath__51__48__I0 (.Y(inst_cellmath__51__48__out0[0]), .A(inst_cellmath__51__48__in1[8]), .B(inst_cellmath__51__48__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__51_0_bdw2052368036_bdw (
	inst_cellmath__51_0_out0,
	inst_cellmath__51_0_in0,
	inst_cellmath__51_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__51_0_out0;
input [0:0] inst_cellmath__51_0_in0;
input [9:9] inst_cellmath__51_0_in1;
NOR2BX1 inst_cellmath__51_0_I3 (.Y(inst_cellmath__51_0_out0), .AN(inst_cellmath__51_0_in0[0]), .B(inst_cellmath__51_0_in1[9]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__28_0_bdw2052368036_bdw (
	inst_cellmath__28_0_out0,
	inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__28_0_out0;
input  inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1;
OR2XL inst_cellmath__28_0_I0 (.Y(inst_cellmath__28_0_out0), .A(inst_cellmath__28_0_in0), .B(inst_cellmath__28_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__27_0_bdw2052368036_bdw (
	inst_cellmath__27_0_out0,
	inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__27_0_out0;
input  inst_cellmath__27_0_in0,
	inst_cellmath__27_0_in1;
OR2XL inst_cellmath__27_0_I0 (.Y(inst_cellmath__27_0_out0), .A(inst_cellmath__27_0_in0), .B(inst_cellmath__27_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__50__50__bdw2052368036_bdw (
	inst_cellmath__50__50__out0,
	inst_cellmath__50__50__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__50__50__out0;
input [9:0] inst_cellmath__50__50__in0;
wire N13,N14,N18,N21,N22;
NOR2XL inst_cellmath__50__50__I0 (.Y(N13), .A(inst_cellmath__50__50__in0[8]), .B(inst_cellmath__50__50__in0[1]));
NOR2XL inst_cellmath__50__50__I1 (.Y(N14), .A(inst_cellmath__50__50__in0[6]), .B(inst_cellmath__50__50__in0[9]));
NAND2XL inst_cellmath__50__50__I5 (.Y(N18), .A(N13), .B(N14));
NOR4X1 inst_cellmath__50__50__I13 (.Y(N22), .A(inst_cellmath__50__50__in0[0]), .B(inst_cellmath__50__50__in0[2]), .C(inst_cellmath__50__50__in0[4]), .D(inst_cellmath__50__50__in0[5]));
NOR3XL inst_cellmath__50__50__I12 (.Y(N21), .A(inst_cellmath__50__50__in0[7]), .B(inst_cellmath__50__50__in0[3]), .C(N18));
NAND2XL inst_cellmath__50__50__I10 (.Y(inst_cellmath__50__50__out0[0]), .A(N22), .B(N21));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__49_1_bdw2052368036_bdw (
	inst_cellmath__49_1_out0,
	inst_cellmath__49_1_in0,
	inst_cellmath__49_1_in1,
	inst_cellmath__49_1_in2,
	inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5
	); /* architecture "gate_level" */ 
output  inst_cellmath__49_1_out0;
input  inst_cellmath__49_1_in0;
input [0:0] inst_cellmath__49_1_in1;
input [9:9] inst_cellmath__49_1_in2;
input  inst_cellmath__49_1_in3,
	inst_cellmath__49_1_in4,
	inst_cellmath__49_1_in5;
wire N13,N14;
NOR4XL inst_cellmath__49_1_I9 (.Y(N13), .A(inst_cellmath__49_1_in3), .B(inst_cellmath__49_1_in4), .C(inst_cellmath__49_1_in5), .D(inst_cellmath__49_1_in2[9]));
NAND2XL inst_cellmath__49_1_I5 (.Y(N14), .A(N13), .B(inst_cellmath__49_1_in1[0]));
OR2XL inst_cellmath__49_1_I6 (.Y(inst_cellmath__49_1_out0), .A(N14), .B(inst_cellmath__49_1_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__43__bdw2052368036_bdw (
	inst_cellmath__37__43__out0,
	inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__43__out0;
input  inst_cellmath__37__43__in0,
	inst_cellmath__37__43__in1;
OR2XL inst_cellmath__37__43__I0 (.Y(inst_cellmath__37__43__out0[0]), .A(inst_cellmath__37__43__in0), .B(inst_cellmath__37__43__in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__11__bdw2052368036_bdw (
	inst_cellmath__32__11__out0,
	inst_cellmath__32__11__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__32__11__out0;
input [8:7] inst_cellmath__32__11__in0;
OR2XL inst_cellmath__32__11__I0 (.Y(inst_cellmath__32__11__out0[0]), .A(inst_cellmath__32__11__in0[8]), .B(inst_cellmath__32__11__in0[7]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__32__10__bdw2052368036_bdw (
	inst_cellmath__32__10__out0,
	inst_cellmath__32__10__in0,
	inst_cellmath__32__10__in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__32__10__out0;
input [0:0] inst_cellmath__32__10__in0;
input [9:9] inst_cellmath__32__10__in1;
NAND2BXL inst_cellmath__32__10__I2 (.Y(inst_cellmath__32__10__out0), .AN(inst_cellmath__32__10__in1[9]), .B(inst_cellmath__32__10__in0[0]));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__37__42__bdw2052368036_bdw (
	inst_cellmath__37__42__out0,
	inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__37__42__out0;
input  inst_cellmath__37__42__in0,
	inst_cellmath__37__42__in1;
OR2XL inst_cellmath__37__42__I0 (.Y(inst_cellmath__37__42__out0[0]), .A(inst_cellmath__37__42__in1), .B(inst_cellmath__37__42__in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__7_0_bdw2052368036_bdw (
	inst_cellmath__7_0_out0,
	inst_cellmath__7_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__7_0_out0;
input [2:0] inst_cellmath__7_0_in0;
wire N42;
NAND2XL inst_cellmath__7_0_I24 (.Y(N42), .A(inst_cellmath__7_0_in0[0]), .B(inst_cellmath__7_0_in0[1]));
NOR2XL inst_cellmath__7_0_I25 (.Y(inst_cellmath__7_0_out0), .A(inst_cellmath__7_0_in0[2]), .B(N42));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__42_0_bdw2052368036_bdw (
	inst_cellmath__42_0_out0,
	inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3
	); /* architecture "gate_level" */ 
output  inst_cellmath__42_0_out0;
input  inst_cellmath__42_0_in0,
	inst_cellmath__42_0_in1,
	inst_cellmath__42_0_in2,
	inst_cellmath__42_0_in3;
wire N12,N21;
INVXL inst_cellmath__42_0_I6 (.Y(N21), .A(inst_cellmath__42_0_in3));
MXI2XL inst_cellmath__42_0_I3 (.Y(N12), .A(inst_cellmath__42_0_in0), .B(N21), .S0(inst_cellmath__42_0_in1));
MX2XL inst_cellmath__42_0_I4 (.Y(inst_cellmath__42_0_out0), .A(N12), .B(N21), .S0(inst_cellmath__42_0_in2));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__52_0_bdw2052368036_bdw (
	inst_cellmath__52_0_out0,
	inst_cellmath__52_0_in0,
	inst_cellmath__52_0_in1,
	inst_cellmath__52_0_in2,
	inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__52_0_out0;
input  inst_cellmath__52_0_in0;
input [7:0] inst_cellmath__52_0_in1;
input  inst_cellmath__52_0_in2;
input [0:0] inst_cellmath__52_0_in3,
	inst_cellmath__52_0_in4;
wire N50,N134,N137,N138;
INVXL inst_cellmath__52_0_I54 (.Y(N137), .A(inst_cellmath__52_0_in4[0]));
AOI21XL inst_cellmath__52_0_I56 (.Y(N50), .A0(inst_cellmath__52_0_in2), .A1(N137), .B0(inst_cellmath__52_0_in3[0]));
OR2XL inst_cellmath__52_0_I57 (.Y(N134), .A(N137), .B(inst_cellmath__52_0_in3[0]));
INVXL inst_cellmath__52_0_I55 (.Y(N138), .A(inst_cellmath__52_0_in1[0]));
MXI2XL inst_cellmath__52_0_I32 (.Y(inst_cellmath__52_0_out0[0]), .A(N138), .B(N50), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I33 (.Y(inst_cellmath__52_0_out0[1]), .A(inst_cellmath__52_0_in1[1]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I34 (.Y(inst_cellmath__52_0_out0[2]), .A(inst_cellmath__52_0_in1[2]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I35 (.Y(inst_cellmath__52_0_out0[3]), .A(inst_cellmath__52_0_in1[3]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I36 (.Y(inst_cellmath__52_0_out0[4]), .A(inst_cellmath__52_0_in1[4]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I37 (.Y(inst_cellmath__52_0_out0[5]), .A(inst_cellmath__52_0_in1[5]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I38 (.Y(inst_cellmath__52_0_out0[6]), .A(inst_cellmath__52_0_in1[6]), .B(N134), .S0(inst_cellmath__52_0_in0));
MX2XL inst_cellmath__52_0_I39 (.Y(inst_cellmath__52_0_out0[7]), .A(inst_cellmath__52_0_in1[7]), .B(N134), .S0(inst_cellmath__52_0_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__47_0_bdw2052368036_bdw (
	inst_cellmath__47_0_out0,
	inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4
	); /* architecture "gate_level" */ 
output  inst_cellmath__47_0_out0;
input  inst_cellmath__47_0_in0,
	inst_cellmath__47_0_in1,
	inst_cellmath__47_0_in2,
	inst_cellmath__47_0_in3,
	inst_cellmath__47_0_in4;
wire N12;
OR4X1 inst_cellmath__47_0_I7 (.Y(N12), .A(inst_cellmath__47_0_in2), .B(inst_cellmath__47_0_in3), .C(inst_cellmath__47_0_in4), .D(inst_cellmath__47_0_in0));
NOR2XL inst_cellmath__47_0_I5 (.Y(inst_cellmath__47_0_out0), .A(N12), .B(inst_cellmath__47_0_in1));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_U_bdw2052368036_bdw (
	inst_cellmath__53_U_out0,
	inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1,
	inst_cellmath__53_U_in2,
	inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4,
	inst_cellmath__53_U_in5
	); /* architecture "gate_level" */ 
output [22:22] inst_cellmath__53_U_out0;
input  inst_cellmath__53_U_in0,
	inst_cellmath__53_U_in1;
input [22:22] inst_cellmath__53_U_in2;
input  inst_cellmath__53_U_in3,
	inst_cellmath__53_U_in4;
input [46:46] inst_cellmath__53_U_in5;
wire N13,N17;
NOR2XL inst_cellmath__53_U_I1 (.Y(N13), .A(inst_cellmath__53_U_in4), .B(inst_cellmath__53_U_in1));
MXI2XL inst_cellmath__53_U_I6 (.Y(N17), .A(inst_cellmath__53_U_in5[46]), .B(inst_cellmath__53_U_in2[22]), .S0(inst_cellmath__53_U_in3));
MXI2XL inst_cellmath__53_U_I7 (.Y(inst_cellmath__53_U_out0[22]), .A(N17), .B(N13), .S0(inst_cellmath__53_U_in0));
endmodule

module cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2052368036_bdw (
	inst_cellmath__53_M_out0,
	inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1,
	inst_cellmath__53_M_in2,
	inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4,
	inst_cellmath__53_M_in5,
	inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7,
	inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9
	); /* architecture "gate_level" */ 
output [21:0] inst_cellmath__53_M_out0;
input  inst_cellmath__53_M_in0,
	inst_cellmath__53_M_in1;
input [21:0] inst_cellmath__53_M_in2;
input  inst_cellmath__53_M_in3,
	inst_cellmath__53_M_in4;
input [45:24] inst_cellmath__53_M_in5;
input  inst_cellmath__53_M_in6,
	inst_cellmath__53_M_in7;
input [21:0] inst_cellmath__53_M_in8,
	inst_cellmath__53_M_in9;
wire N135,N137,N142,N144,N146,N148,N150 
	,N152,N154,N156,N158,N160,N162,N164,N166 
	,N168,N170,N172,N174,N176,N178,N180,N182 
	,N184,N236,N238,N240,N242,N244,N246,N248 
	,N250,N252,N254,N256,N258,N260,N262,N264 
	,N266,N268,N270,N272,N274,N276,N278,N281 
	,N285,N289,N293,N297,N301,N305,N309,N313 
	,N317,N321,N325,N329,N333,N337,N341,N345 
	,N349,N353,N357,N361,N365,N368,N370,N372 
	,N538,N547,N548;
INVXL inst_cellmath__53_M_I182 (.Y(N538), .A(inst_cellmath__53_M_in0));
NOR2XL inst_cellmath__53_M_I7 (.Y(N368), .A(inst_cellmath__53_M_in4), .B(N538));
NAND3BXL inst_cellmath__53_M_I429 (.Y(N135), .AN(inst_cellmath__53_M_in7), .B(inst_cellmath__53_M_in6), .C(inst_cellmath__53_M_in4));
NOR2XL inst_cellmath__53_M_I11 (.Y(N370), .A(N135), .B(N538));
NAND2XL inst_cellmath__53_M_I12 (.Y(N137), .A(inst_cellmath__53_M_in7), .B(inst_cellmath__53_M_in4));
NOR2XL inst_cellmath__53_M_I13 (.Y(N372), .A(N137), .B(N538));
NOR2BX1 inst_cellmath__53_M_I200 (.Y(N547), .AN(N538), .B(inst_cellmath__53_M_in3));
AND2XL inst_cellmath__53_M_I201 (.Y(N548), .A(inst_cellmath__53_M_in3), .B(N538));
AOI22XL inst_cellmath__53_M_I17 (.Y(N142), .A0(inst_cellmath__53_M_in2[0]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[24]));
AOI22XL inst_cellmath__53_M_I18 (.Y(N144), .A0(inst_cellmath__53_M_in2[1]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[25]));
AOI22XL inst_cellmath__53_M_I19 (.Y(N146), .A0(inst_cellmath__53_M_in2[2]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[26]));
AOI22XL inst_cellmath__53_M_I20 (.Y(N148), .A0(inst_cellmath__53_M_in2[3]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[27]));
AOI22XL inst_cellmath__53_M_I21 (.Y(N150), .A0(inst_cellmath__53_M_in2[4]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[28]));
AOI22XL inst_cellmath__53_M_I22 (.Y(N152), .A0(inst_cellmath__53_M_in2[5]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[29]));
AOI22XL inst_cellmath__53_M_I23 (.Y(N154), .A0(inst_cellmath__53_M_in2[6]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[30]));
AOI22XL inst_cellmath__53_M_I24 (.Y(N156), .A0(inst_cellmath__53_M_in2[7]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[31]));
AOI22XL inst_cellmath__53_M_I25 (.Y(N158), .A0(inst_cellmath__53_M_in2[8]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[32]));
AOI22XL inst_cellmath__53_M_I26 (.Y(N160), .A0(inst_cellmath__53_M_in2[9]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[33]));
AOI22XL inst_cellmath__53_M_I27 (.Y(N162), .A0(inst_cellmath__53_M_in2[10]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[34]));
AOI22XL inst_cellmath__53_M_I28 (.Y(N164), .A0(inst_cellmath__53_M_in2[11]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[35]));
AOI22XL inst_cellmath__53_M_I29 (.Y(N166), .A0(inst_cellmath__53_M_in2[12]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[36]));
AOI22XL inst_cellmath__53_M_I30 (.Y(N168), .A0(inst_cellmath__53_M_in2[13]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[37]));
AOI22XL inst_cellmath__53_M_I31 (.Y(N170), .A0(inst_cellmath__53_M_in2[14]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[38]));
AOI22XL inst_cellmath__53_M_I32 (.Y(N172), .A0(inst_cellmath__53_M_in2[15]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[39]));
AOI22XL inst_cellmath__53_M_I33 (.Y(N174), .A0(inst_cellmath__53_M_in2[16]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[40]));
AOI22XL inst_cellmath__53_M_I34 (.Y(N176), .A0(inst_cellmath__53_M_in2[17]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[41]));
AOI22XL inst_cellmath__53_M_I35 (.Y(N178), .A0(inst_cellmath__53_M_in2[18]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[42]));
AOI22XL inst_cellmath__53_M_I36 (.Y(N180), .A0(inst_cellmath__53_M_in2[19]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[43]));
AOI22XL inst_cellmath__53_M_I37 (.Y(N182), .A0(inst_cellmath__53_M_in2[20]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[44]));
AOI22XL inst_cellmath__53_M_I38 (.Y(N184), .A0(inst_cellmath__53_M_in2[21]), .A1(N548), .B0(N547), .B1(inst_cellmath__53_M_in5[45]));
AOI22XL inst_cellmath__53_M_I42 (.Y(N281), .A0(inst_cellmath__53_M_in8[0]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I43 (.Y(N285), .A0(inst_cellmath__53_M_in8[1]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I44 (.Y(N289), .A0(inst_cellmath__53_M_in8[2]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I45 (.Y(N293), .A0(inst_cellmath__53_M_in8[3]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I46 (.Y(N297), .A0(inst_cellmath__53_M_in8[4]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I47 (.Y(N301), .A0(inst_cellmath__53_M_in8[5]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I48 (.Y(N305), .A0(inst_cellmath__53_M_in8[6]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I49 (.Y(N309), .A0(inst_cellmath__53_M_in8[7]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I50 (.Y(N313), .A0(inst_cellmath__53_M_in8[8]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I51 (.Y(N317), .A0(inst_cellmath__53_M_in8[9]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I52 (.Y(N321), .A0(inst_cellmath__53_M_in8[10]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I53 (.Y(N325), .A0(inst_cellmath__53_M_in8[11]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I54 (.Y(N329), .A0(inst_cellmath__53_M_in8[12]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I55 (.Y(N333), .A0(inst_cellmath__53_M_in8[13]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I56 (.Y(N337), .A0(inst_cellmath__53_M_in8[14]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I57 (.Y(N341), .A0(inst_cellmath__53_M_in8[15]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I58 (.Y(N345), .A0(inst_cellmath__53_M_in8[16]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I59 (.Y(N349), .A0(inst_cellmath__53_M_in8[17]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I60 (.Y(N353), .A0(inst_cellmath__53_M_in8[18]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I61 (.Y(N357), .A0(inst_cellmath__53_M_in8[19]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I62 (.Y(N361), .A0(inst_cellmath__53_M_in8[20]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
AOI22XL inst_cellmath__53_M_I63 (.Y(N365), .A0(inst_cellmath__53_M_in8[21]), .A1(N370), .B0(N368), .B1(inst_cellmath__53_M_in1));
NAND2XL inst_cellmath__53_M_I67 (.Y(N236), .A(N372), .B(inst_cellmath__53_M_in9[0]));
NAND2XL inst_cellmath__53_M_I68 (.Y(N238), .A(N372), .B(inst_cellmath__53_M_in9[1]));
NAND2XL inst_cellmath__53_M_I69 (.Y(N240), .A(N372), .B(inst_cellmath__53_M_in9[2]));
NAND2XL inst_cellmath__53_M_I70 (.Y(N242), .A(N372), .B(inst_cellmath__53_M_in9[3]));
NAND2XL inst_cellmath__53_M_I71 (.Y(N244), .A(N372), .B(inst_cellmath__53_M_in9[4]));
NAND2XL inst_cellmath__53_M_I72 (.Y(N246), .A(N372), .B(inst_cellmath__53_M_in9[5]));
NAND2XL inst_cellmath__53_M_I73 (.Y(N248), .A(N372), .B(inst_cellmath__53_M_in9[6]));
NAND2XL inst_cellmath__53_M_I74 (.Y(N250), .A(N372), .B(inst_cellmath__53_M_in9[7]));
NAND2XL inst_cellmath__53_M_I75 (.Y(N252), .A(N372), .B(inst_cellmath__53_M_in9[8]));
NAND2XL inst_cellmath__53_M_I76 (.Y(N254), .A(N372), .B(inst_cellmath__53_M_in9[9]));
NAND2XL inst_cellmath__53_M_I77 (.Y(N256), .A(N372), .B(inst_cellmath__53_M_in9[10]));
NAND2XL inst_cellmath__53_M_I78 (.Y(N258), .A(N372), .B(inst_cellmath__53_M_in9[11]));
NAND2XL inst_cellmath__53_M_I79 (.Y(N260), .A(N372), .B(inst_cellmath__53_M_in9[12]));
NAND2XL inst_cellmath__53_M_I80 (.Y(N262), .A(N372), .B(inst_cellmath__53_M_in9[13]));
NAND2XL inst_cellmath__53_M_I81 (.Y(N264), .A(N372), .B(inst_cellmath__53_M_in9[14]));
NAND2XL inst_cellmath__53_M_I82 (.Y(N266), .A(N372), .B(inst_cellmath__53_M_in9[15]));
NAND2XL inst_cellmath__53_M_I83 (.Y(N268), .A(N372), .B(inst_cellmath__53_M_in9[16]));
NAND2XL inst_cellmath__53_M_I84 (.Y(N270), .A(N372), .B(inst_cellmath__53_M_in9[17]));
NAND2XL inst_cellmath__53_M_I85 (.Y(N272), .A(N372), .B(inst_cellmath__53_M_in9[18]));
NAND2XL inst_cellmath__53_M_I86 (.Y(N274), .A(N372), .B(inst_cellmath__53_M_in9[19]));
NAND2XL inst_cellmath__53_M_I87 (.Y(N276), .A(N372), .B(inst_cellmath__53_M_in9[20]));
NAND2XL inst_cellmath__53_M_I88 (.Y(N278), .A(N372), .B(inst_cellmath__53_M_in9[21]));
NAND3XL inst_cellmath__53_M_I202 (.Y(inst_cellmath__53_M_out0[0]), .A(N236), .B(N142), .C(N281));
NAND3XL inst_cellmath__53_M_I203 (.Y(inst_cellmath__53_M_out0[1]), .A(N238), .B(N144), .C(N285));
NAND3XL inst_cellmath__53_M_I204 (.Y(inst_cellmath__53_M_out0[2]), .A(N240), .B(N146), .C(N289));
NAND3XL inst_cellmath__53_M_I205 (.Y(inst_cellmath__53_M_out0[3]), .A(N242), .B(N148), .C(N293));
NAND3XL inst_cellmath__53_M_I206 (.Y(inst_cellmath__53_M_out0[4]), .A(N244), .B(N150), .C(N297));
NAND3XL inst_cellmath__53_M_I207 (.Y(inst_cellmath__53_M_out0[5]), .A(N246), .B(N152), .C(N301));
NAND3XL inst_cellmath__53_M_I208 (.Y(inst_cellmath__53_M_out0[6]), .A(N248), .B(N154), .C(N305));
NAND3XL inst_cellmath__53_M_I209 (.Y(inst_cellmath__53_M_out0[7]), .A(N250), .B(N156), .C(N309));
NAND3XL inst_cellmath__53_M_I210 (.Y(inst_cellmath__53_M_out0[8]), .A(N252), .B(N158), .C(N313));
NAND3XL inst_cellmath__53_M_I211 (.Y(inst_cellmath__53_M_out0[9]), .A(N254), .B(N160), .C(N317));
NAND3XL inst_cellmath__53_M_I212 (.Y(inst_cellmath__53_M_out0[10]), .A(N256), .B(N162), .C(N321));
NAND3XL inst_cellmath__53_M_I213 (.Y(inst_cellmath__53_M_out0[11]), .A(N258), .B(N164), .C(N325));
NAND3XL inst_cellmath__53_M_I214 (.Y(inst_cellmath__53_M_out0[12]), .A(N260), .B(N166), .C(N329));
NAND3XL inst_cellmath__53_M_I215 (.Y(inst_cellmath__53_M_out0[13]), .A(N262), .B(N168), .C(N333));
NAND3XL inst_cellmath__53_M_I216 (.Y(inst_cellmath__53_M_out0[14]), .A(N264), .B(N170), .C(N337));
NAND3XL inst_cellmath__53_M_I217 (.Y(inst_cellmath__53_M_out0[15]), .A(N266), .B(N172), .C(N341));
NAND3XL inst_cellmath__53_M_I218 (.Y(inst_cellmath__53_M_out0[16]), .A(N268), .B(N174), .C(N345));
NAND3XL inst_cellmath__53_M_I219 (.Y(inst_cellmath__53_M_out0[17]), .A(N270), .B(N176), .C(N349));
NAND3XL inst_cellmath__53_M_I220 (.Y(inst_cellmath__53_M_out0[18]), .A(N272), .B(N178), .C(N353));
NAND3XL inst_cellmath__53_M_I221 (.Y(inst_cellmath__53_M_out0[19]), .A(N274), .B(N180), .C(N357));
NAND3XL inst_cellmath__53_M_I222 (.Y(inst_cellmath__53_M_out0[20]), .A(N276), .B(N182), .C(N361));
NAND3XL inst_cellmath__53_M_I223 (.Y(inst_cellmath__53_M_out0[21]), .A(N278), .B(N184), .C(N365));
endmodule

/* CADENCE  ubLxSQzXqR0= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/




module float_div_cynw_cm_float_mul_ieee_E8_M23_5( a_sign, a_exp, a_man, b_sign, b_exp, b_man, rm, x, aclk, astall );
input a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire[31:0] x_wire;
input aclk;
input astall;
cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2052368036_bdw cynw_cm_float_mul_ieee_inst_cellmath__53_M_bdw2469856145_bdw_inst( .a_sign(a_sign), .a_exp(a_exp), .a_man(a_man), .b_sign(b_sign), .b_exp(b_exp), .b_man(b_man), .rm(rm), .x(x_wire));
reg [31:0] x_reg_0;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_0 <= x_wire;
end
/* $A : movable_reg = reset */
reg [31:0] x_reg_1;
/* $A : movable_reg */
always @(posedge aclk) begin
    if ( !astall) x_reg_1 <= x_reg_0;
end
/* $A : movable_reg = reset */
assign x = x_reg_1;
endmodule


