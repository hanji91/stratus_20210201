/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:05 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_5 (
	a_sign,
	a_exp,
	a_man,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [36:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_x;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19;
wire [7:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20;
wire [8:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42;
wire [18:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51;
wire [24:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60;
wire [39:0] float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64;
wire  float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743,
	float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
wire N5677,N5682,N5687,N5692,N5697,N5702,N5707 
	,N5712,N5717,N11884,N11888,N11890,N12051,N12056,N12061 
	,N12066,N12071,N12076,N12164,N12168,N12170,N12229,N12234 
	,N12239,N12244,N12249,N12254,N12259,N12266,N12274,N12291 
	,N12295,N12309,N12317,N12325,N12333,N12349,N12365,N12416 
	,N12418,N12420,N12445,N12449,N12511,N12513,N12546,N12581 
	,N12587,N12589,N12622,N12628,N12663,N12704,N12724,N12726 
	,N12728,N12769,N12777,N12781,N12822,N12881,N12895,N12945 
	,N12967,N12975,N12977,N12979,N13040,N13048,N13060,N13066 
	,N13068,N13070,N13129,N13145,N13153,N13155,N13157,N13215 
	,N13223,N13235,N13241,N13243,N13245,N13254,N13261,N13263 
	,N13319,N13364,N13366,N13432,N13455,N13465,N13470,N13476 
	,N13478,N13494,N13496,N13498,N13610,N13616,N13618,N13624 
	,N13626,N13628,N13706,N13712,N13720,N13727,N13735,N13745 
	,N13751,N13753,N13755,N13759,N13761,N13767,N13769,N13771 
	,N13780,N13782,N13784,N13849,N13859,N13867,N13869,N13883 
	,N13885,N13889,N13907,N13917,N13925,N13931,N13933,N13935 
	,N13944,N13946,N13948,N14002,N14006,N14014,N14018,N14024 
	,N14030,N14038,N14040,N14060,N14071,N14073,N14075,N14079 
	,N14081,N14083,N14087,N14089,N14091,N14158,N14160,N14166 
	,N14168,N14174,N14178,N14182,N14184,N14186,N14202,N14204 
	,N14206,N14209,N14214,N14230,N14232,N14234,N14260,N14278 
	,N14284,N14286,N14288,N14292,N14294,N14296,N14301,N14316 
	,N14318,N14320,N14324,N14326,N14328,N14339,N14370,N14374 
	,N14376,N14378,N14382,N14384,N14386,N14390,N14392,N14394 
	,N14398,N14400,N14402,N14406,N14408,N14419,N14421,N14423 
	,N14435,N14441,N14443,N14454,N14456,N14465,N14469,N14471 
	,N14473,N14479,N14481,N14483,N14487,N14489,N14491,N14494 
	,N14505,N14507,N14509,N14515,N14517,N14519,N14526,N14535 
	,N14543,N14551,N14556,N14562,N15230,N15238,N15245,N15271 
	,N15281,N15285,N15287,N15289,N15293,N15832,N15834,N15845 
	,N15848,N15849,N15851,N15853,N15854,N15856,N15858,N15860 
	,N15861,N15863,N15865,N15867,N15869,N15870,N15871,N15873 
	,N15875,N15878,N15881,N15883,N15885,N15886,N15888,N15894 
	,N15929,N15933,N15934,N15935,N15936,N15939,N15940,N15942 
	,N15944,N15947,N15949,N15952,N15957,N15959,N15963,N15993 
	,N15996,N15997,N16001,N16003,N16005,N16008,N16010,N16012 
	,N16014,N16016,N16017,N16019,N16020,N16022,N16025,N16027 
	,N16029,N16030,N16032,N16034,N16038,N16039,N16040,N16042 
	,N16075,N16079,N16080,N16082,N16084,N16085,N16087,N16089 
	,N16091,N16093,N16095,N16099,N16101,N16102,N16104,N16105 
	,N16107,N16108,N16111,N16113,N16115,N16116,N16119,N16120 
	,N16121,N16123,N16126,N16128,N16162,N16165,N16167,N16168 
	,N16169,N16171,N16173,N16185,N16186,N16190,N16193,N16194 
	,N16197,N16199,N16201,N16203;
reg x_reg_L1_22__retimed_I8255_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I8255_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736;
	end
assign N15293 = x_reg_L1_22__retimed_I8255_QOUT;
reg x_reg_L1_22__retimed_I8254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I8254_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13];
	end
assign x[13] = x_reg_L1_22__retimed_I8254_QOUT;
reg x_reg_L0_22__retimed_I8253_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8253_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919;
	end
assign N15289 = x_reg_L0_22__retimed_I8253_QOUT;
reg x_reg_L0_22__retimed_I8252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8252_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409;
	end
assign N15287 = x_reg_L0_22__retimed_I8252_QOUT;
reg x_reg_L0_22__retimed_I8251_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8251_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777;
	end
assign N15285 = x_reg_L0_22__retimed_I8251_QOUT;
reg x_reg_L0_22__retimed_I8250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8250_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305;
	end
assign N15281 = x_reg_L0_22__retimed_I8250_QOUT;
reg x_reg_L0_22__retimed_I8246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8246_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803;
	end
assign N15271 = x_reg_L0_22__retimed_I8246_QOUT;
reg x_reg_L0_22__retimed_I8235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8235_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294;
	end
assign N15245 = x_reg_L0_22__retimed_I8235_QOUT;
reg x_reg_L0_22__retimed_I8232_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8232_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134;
	end
assign N15238 = x_reg_L0_22__retimed_I8232_QOUT;
reg x_reg_L0_22__retimed_I8229_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I8229_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221;
	end
assign N15230 = x_reg_L0_22__retimed_I8229_QOUT;
reg x_reg_L0_22__retimed_I7935_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7935_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640;
	end
assign N14519 = x_reg_L0_22__retimed_I7935_QOUT;
reg x_reg_L0_22__retimed_I7934_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7934_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884;
	end
assign N14517 = x_reg_L0_22__retimed_I7934_QOUT;
reg x_reg_L0_22__retimed_I7933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7933_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5];
	end
assign N14515 = x_reg_L0_22__retimed_I7933_QOUT;
reg x_reg_L0_22__retimed_I7932_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7932_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212;
	end
assign N14509 = x_reg_L0_22__retimed_I7932_QOUT;
reg x_reg_L0_22__retimed_I7931_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7931_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839;
	end
assign N14507 = x_reg_L0_22__retimed_I7931_QOUT;
reg x_reg_L0_22__retimed_I7930_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7930_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357;
	end
assign N14505 = x_reg_L0_22__retimed_I7930_QOUT;
reg x_reg_L0_22__retimed_I7926_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7926_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748;
	end
assign N14494 = x_reg_L0_22__retimed_I7926_QOUT;
reg x_reg_L0_22__retimed_I7925_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7925_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7];
	end
assign N14491 = x_reg_L0_22__retimed_I7925_QOUT;
reg x_reg_L0_22__retimed_I7924_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7924_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7];
	end
assign N14489 = x_reg_L0_22__retimed_I7924_QOUT;
reg x_reg_L0_22__retimed_I7923_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7923_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7];
	end
assign N14487 = x_reg_L0_22__retimed_I7923_QOUT;
reg x_reg_L0_22__retimed_I7922_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7922_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542;
	end
assign N14483 = x_reg_L0_22__retimed_I7922_QOUT;
reg x_reg_L0_22__retimed_I7921_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7921_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667;
	end
assign N14481 = x_reg_L0_22__retimed_I7921_QOUT;
reg x_reg_L0_22__retimed_I7920_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7920_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6];
	end
assign N14479 = x_reg_L0_22__retimed_I7920_QOUT;
reg x_reg_L0_22__retimed_I7919_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7919_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772;
	end
assign N14473 = x_reg_L0_22__retimed_I7919_QOUT;
reg x_reg_L0_22__retimed_I7918_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7918_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255;
	end
assign N14471 = x_reg_L0_22__retimed_I7918_QOUT;
reg x_reg_L0_22__retimed_I7917_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7917_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404;
	end
assign N14469 = x_reg_L0_22__retimed_I7917_QOUT;
reg x_reg_L0_22__retimed_I7916_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7916_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605;
	end
assign N14465 = x_reg_L0_22__retimed_I7916_QOUT;
reg x_reg_L0_22__retimed_I7912_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7912_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8];
	end
assign N14456 = x_reg_L0_22__retimed_I7912_QOUT;
reg x_reg_L0_22__retimed_I7911_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7911_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8];
	end
assign N14454 = x_reg_L0_22__retimed_I7911_QOUT;
reg x_reg_L0_22__retimed_I7907_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7907_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451;
	end
assign N14443 = x_reg_L0_22__retimed_I7907_QOUT;
reg x_reg_L0_22__retimed_I7906_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7906_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7];
	end
assign N14441 = x_reg_L0_22__retimed_I7906_QOUT;
reg x_reg_L0_22__retimed_I7905_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7905_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22];
	end
assign N14435 = x_reg_L0_22__retimed_I7905_QOUT;
reg x_reg_L0_22__retimed_I7904_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7904_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194;
	end
assign N14423 = x_reg_L0_22__retimed_I7904_QOUT;
reg x_reg_L0_22__retimed_I7903_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7903_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069;
	end
assign N14421 = x_reg_L0_22__retimed_I7903_QOUT;
reg x_reg_L0_22__retimed_I7902_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7902_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201;
	end
assign N14419 = x_reg_L0_22__retimed_I7902_QOUT;
reg x_reg_L0_22__retimed_I7898_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7898_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769;
	end
assign N14408 = x_reg_L0_22__retimed_I7898_QOUT;
reg x_reg_L0_22__retimed_I7897_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7897_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811;
	end
assign N14406 = x_reg_L0_22__retimed_I7897_QOUT;
reg x_reg_L0_22__retimed_I7896_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7896_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216;
	end
assign N14402 = x_reg_L0_22__retimed_I7896_QOUT;
reg x_reg_L0_22__retimed_I7895_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7895_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282;
	end
assign N14400 = x_reg_L0_22__retimed_I7895_QOUT;
reg x_reg_L0_22__retimed_I7894_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7894_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078;
	end
assign N14398 = x_reg_L0_22__retimed_I7894_QOUT;
reg x_reg_L0_22__retimed_I7893_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7893_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571;
	end
assign N14394 = x_reg_L0_22__retimed_I7893_QOUT;
reg x_reg_L0_22__retimed_I7892_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7892_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960;
	end
assign N14392 = x_reg_L0_22__retimed_I7892_QOUT;
reg x_reg_L0_22__retimed_I7891_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7891_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195;
	end
assign N14390 = x_reg_L0_22__retimed_I7891_QOUT;
reg x_reg_L0_22__retimed_I7890_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7890_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180;
	end
assign N14386 = x_reg_L0_22__retimed_I7890_QOUT;
reg x_reg_L0_22__retimed_I7889_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7889_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340;
	end
assign N14384 = x_reg_L0_22__retimed_I7889_QOUT;
reg x_reg_L0_22__retimed_I7888_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7888_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373;
	end
assign N14382 = x_reg_L0_22__retimed_I7888_QOUT;
reg x_reg_L0_22__retimed_I7887_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7887_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077;
	end
assign N14378 = x_reg_L0_22__retimed_I7887_QOUT;
reg x_reg_L0_22__retimed_I7886_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7886_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266;
	end
assign N14376 = x_reg_L0_22__retimed_I7886_QOUT;
reg x_reg_L0_22__retimed_I7885_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7885_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235;
	end
assign N14374 = x_reg_L0_22__retimed_I7885_QOUT;
reg x_reg_L0_22__retimed_I7884_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7884_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9];
	end
assign N14370 = x_reg_L0_22__retimed_I7884_QOUT;
reg x_reg_L0_22__retimed_I7871_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7871_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8];
	end
assign N14339 = x_reg_L0_22__retimed_I7871_QOUT;
reg x_reg_L0_22__retimed_I7868_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7868_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252;
	end
assign N14328 = x_reg_L0_22__retimed_I7868_QOUT;
reg x_reg_L0_22__retimed_I7867_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7867_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093;
	end
assign N14326 = x_reg_L0_22__retimed_I7867_QOUT;
reg x_reg_L0_22__retimed_I7866_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7866_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108;
	end
assign N14324 = x_reg_L0_22__retimed_I7866_QOUT;
reg x_reg_L0_22__retimed_I7865_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7865_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304;
	end
assign N14320 = x_reg_L0_22__retimed_I7865_QOUT;
reg x_reg_L0_22__retimed_I7864_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7864_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169;
	end
assign N14318 = x_reg_L0_22__retimed_I7864_QOUT;
reg x_reg_L0_22__retimed_I7863_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7863_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091;
	end
assign N14316 = x_reg_L0_22__retimed_I7863_QOUT;
reg x_reg_L0_22__retimed_I7861_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7861_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588;
	end
assign N14301 = x_reg_L0_22__retimed_I7861_QOUT;
reg x_reg_L0_22__retimed_I7859_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7859_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021;
	end
assign N14296 = x_reg_L0_22__retimed_I7859_QOUT;
reg x_reg_L0_22__retimed_I7858_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7858_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895;
	end
assign N14294 = x_reg_L0_22__retimed_I7858_QOUT;
reg x_reg_L0_22__retimed_I7857_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7857_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508;
	end
assign N14292 = x_reg_L0_22__retimed_I7857_QOUT;
reg x_reg_L0_22__retimed_I7856_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7856_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365;
	end
assign N14288 = x_reg_L0_22__retimed_I7856_QOUT;
reg x_reg_L0_22__retimed_I7855_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7855_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160;
	end
assign N14286 = x_reg_L0_22__retimed_I7855_QOUT;
reg x_reg_L0_22__retimed_I7854_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7854_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293;
	end
assign N14284 = x_reg_L0_22__retimed_I7854_QOUT;
reg x_reg_L0_22__retimed_I7852_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7852_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240;
	end
assign N14278 = x_reg_L0_22__retimed_I7852_QOUT;
reg x_reg_L0_22__retimed_I7845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7845_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153;
	end
assign N14260 = x_reg_L0_22__retimed_I7845_QOUT;
reg x_reg_L0_22__retimed_I7836_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7836_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156;
	end
assign N14234 = x_reg_L0_22__retimed_I7836_QOUT;
reg x_reg_L0_22__retimed_I7835_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7835_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521;
	end
assign N14232 = x_reg_L0_22__retimed_I7835_QOUT;
reg x_reg_L0_22__retimed_I7834_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7834_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784;
	end
assign N14230 = x_reg_L0_22__retimed_I7834_QOUT;
reg x_reg_L0_22__retimed_I7828_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7828_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324;
	end
assign N14214 = x_reg_L0_22__retimed_I7828_QOUT;
reg x_reg_L0_22__retimed_I7826_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7826_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248;
	end
assign N14209 = x_reg_L0_22__retimed_I7826_QOUT;
reg x_reg_L0_22__retimed_I7825_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7825_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238;
	end
assign N14206 = x_reg_L0_22__retimed_I7825_QOUT;
reg x_reg_L0_22__retimed_I7824_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7824_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374;
	end
assign N14204 = x_reg_L0_22__retimed_I7824_QOUT;
reg x_reg_L0_22__retimed_I7823_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7823_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168;
	end
assign N14202 = x_reg_L0_22__retimed_I7823_QOUT;
reg x_reg_L0_22__retimed_I7821_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7821_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846;
	end
assign N14186 = x_reg_L0_22__retimed_I7821_QOUT;
reg x_reg_L0_22__retimed_I7820_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7820_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332;
	end
assign N14184 = x_reg_L0_22__retimed_I7820_QOUT;
reg x_reg_L0_22__retimed_I7819_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7819_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208;
	end
assign N14182 = x_reg_L0_22__retimed_I7819_QOUT;
reg x_reg_L0_22__retimed_I7818_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7818_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114;
	end
assign N14178 = x_reg_L0_22__retimed_I7818_QOUT;
reg x_reg_L0_22__retimed_I7816_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7816_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315;
	end
assign N14174 = x_reg_L0_22__retimed_I7816_QOUT;
reg x_reg_L0_22__retimed_I7814_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7814_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380;
	end
assign N14168 = x_reg_L0_22__retimed_I7814_QOUT;
reg x_reg_L0_22__retimed_I7813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7813_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306;
	end
assign N14166 = x_reg_L0_22__retimed_I7813_QOUT;
reg x_reg_L0_22__retimed_I7811_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7811_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186;
	end
assign N14160 = x_reg_L0_22__retimed_I7811_QOUT;
reg x_reg_L0_22__retimed_I7810_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7810_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322;
	end
assign N14158 = x_reg_L0_22__retimed_I7810_QOUT;
reg x_reg_L0_22__retimed_I7785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7785_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859;
	end
assign N14091 = x_reg_L0_22__retimed_I7785_QOUT;
reg x_reg_L0_22__retimed_I7784_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7784_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872;
	end
assign N14089 = x_reg_L0_22__retimed_I7784_QOUT;
reg x_reg_L0_22__retimed_I7783_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7783_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347;
	end
assign N14087 = x_reg_L0_22__retimed_I7783_QOUT;
reg x_reg_L0_22__retimed_I7782_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7782_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206;
	end
assign N14083 = x_reg_L0_22__retimed_I7782_QOUT;
reg x_reg_L0_22__retimed_I7781_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7781_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200;
	end
assign N14081 = x_reg_L0_22__retimed_I7781_QOUT;
reg x_reg_L0_22__retimed_I7780_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7780_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135;
	end
assign N14079 = x_reg_L0_22__retimed_I7780_QOUT;
reg x_reg_L0_22__retimed_I7779_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7779_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330;
	end
assign N14075 = x_reg_L0_22__retimed_I7779_QOUT;
reg x_reg_L0_22__retimed_I7778_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7778_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124;
	end
assign N14073 = x_reg_L0_22__retimed_I7778_QOUT;
reg x_reg_L0_22__retimed_I7777_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7777_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391;
	end
assign N14071 = x_reg_L0_22__retimed_I7777_QOUT;
reg x_reg_L0_22__retimed_I7773_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7773_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399;
	end
assign N14060 = x_reg_L0_22__retimed_I7773_QOUT;
reg x_reg_L0_22__retimed_I7765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7765_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032;
	end
assign N14040 = x_reg_L0_22__retimed_I7765_QOUT;
reg x_reg_L0_22__retimed_I7764_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7764_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537;
	end
assign N14038 = x_reg_L0_22__retimed_I7764_QOUT;
reg x_reg_L0_22__retimed_I7761_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7761_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116;
	end
assign N14030 = x_reg_L0_22__retimed_I7761_QOUT;
reg x_reg_L0_22__retimed_I7759_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7759_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398;
	end
assign N14024 = x_reg_L0_22__retimed_I7759_QOUT;
reg x_reg_L0_22__retimed_I7757_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7757_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205;
	end
assign N14018 = x_reg_L0_22__retimed_I7757_QOUT;
reg x_reg_L0_22__retimed_I7755_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7755_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397;
	end
assign N14014 = x_reg_L0_22__retimed_I7755_QOUT;
reg x_reg_L0_22__retimed_I7752_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7752_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132;
	end
assign N14006 = x_reg_L0_22__retimed_I7752_QOUT;
reg x_reg_L0_22__retimed_I7751_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7751_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152;
	end
assign N14002 = x_reg_L0_22__retimed_I7751_QOUT;
reg x_reg_L0_22__retimed_I7731_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7731_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532;
	end
assign N13948 = x_reg_L0_22__retimed_I7731_QOUT;
reg x_reg_L0_22__retimed_I7730_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7730_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547;
	end
assign N13946 = x_reg_L0_22__retimed_I7730_QOUT;
reg x_reg_L0_22__retimed_I7729_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7729_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152;
	end
assign N13944 = x_reg_L0_22__retimed_I7729_QOUT;
reg x_reg_L0_22__retimed_I7726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7726_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437;
	end
assign N13935 = x_reg_L0_22__retimed_I7726_QOUT;
reg x_reg_L0_22__retimed_I7725_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7725_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343;
	end
assign N13933 = x_reg_L0_22__retimed_I7725_QOUT;
reg x_reg_L0_22__retimed_I7724_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7724_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967;
	end
assign N13931 = x_reg_L0_22__retimed_I7724_QOUT;
reg x_reg_L0_22__retimed_I7722_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7722_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207;
	end
assign N13925 = x_reg_L0_22__retimed_I7722_QOUT;
reg x_reg_L0_22__retimed_I7719_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7719_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150;
	end
assign N13917 = x_reg_L0_22__retimed_I7719_QOUT;
reg x_reg_L0_22__retimed_I7715_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7715_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248;
	end
assign N13907 = x_reg_L0_22__retimed_I7715_QOUT;
reg x_reg_L0_22__retimed_I7708_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7708_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217;
	end
assign N13889 = x_reg_L0_22__retimed_I7708_QOUT;
reg x_reg_L0_22__retimed_I7707_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7707_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389;
	end
assign N13885 = x_reg_L0_22__retimed_I7707_QOUT;
reg x_reg_L0_22__retimed_I7706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7706_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145;
	end
assign N13883 = x_reg_L0_22__retimed_I7706_QOUT;
reg x_reg_L0_22__retimed_I7701_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7701_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372;
	end
assign N13869 = x_reg_L0_22__retimed_I7701_QOUT;
reg x_reg_L0_22__retimed_I7700_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7700_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225;
	end
assign N13867 = x_reg_L0_22__retimed_I7700_QOUT;
reg x_reg_L0_22__retimed_I7697_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7697_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313;
	end
assign N13859 = x_reg_L0_22__retimed_I7697_QOUT;
reg x_reg_L0_22__retimed_I7693_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7693_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298;
	end
assign N13849 = x_reg_L0_22__retimed_I7693_QOUT;
reg x_reg_L0_22__retimed_I7669_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7669_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147;
	end
assign N13784 = x_reg_L0_22__retimed_I7669_QOUT;
reg x_reg_L0_22__retimed_I7668_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7668_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246;
	end
assign N13782 = x_reg_L0_22__retimed_I7668_QOUT;
reg x_reg_L0_22__retimed_I7667_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7667_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774;
	end
assign N13780 = x_reg_L0_22__retimed_I7667_QOUT;
reg x_reg_L0_22__retimed_I7664_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7664_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435;
	end
assign N13771 = x_reg_L0_22__retimed_I7664_QOUT;
reg x_reg_L0_22__retimed_I7663_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7663_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040;
	end
assign N13769 = x_reg_L0_22__retimed_I7663_QOUT;
reg x_reg_L0_22__retimed_I7662_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7662_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057;
	end
assign N13767 = x_reg_L0_22__retimed_I7662_QOUT;
reg x_reg_L0_22__retimed_I7660_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7660_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527;
	end
assign N13761 = x_reg_L0_22__retimed_I7660_QOUT;
reg x_reg_L0_22__retimed_I7659_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7659_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760;
	end
assign N13759 = x_reg_L0_22__retimed_I7659_QOUT;
reg x_reg_L0_22__retimed_I7658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7658_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297;
	end
assign N13755 = x_reg_L0_22__retimed_I7658_QOUT;
reg x_reg_L0_22__retimed_I7657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7657_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089;
	end
assign N13753 = x_reg_L0_22__retimed_I7657_QOUT;
reg x_reg_L0_22__retimed_I7656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7656_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159;
	end
assign N13751 = x_reg_L0_22__retimed_I7656_QOUT;
reg x_reg_L0_22__retimed_I7654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7654_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280;
	end
assign N13745 = x_reg_L0_22__retimed_I7654_QOUT;
reg x_reg_L0_22__retimed_I7650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7650_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477;
	end
assign N13735 = x_reg_L0_22__retimed_I7650_QOUT;
reg x_reg_L0_22__retimed_I7647_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7647_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855;
	end
assign N13727 = x_reg_L0_22__retimed_I7647_QOUT;
reg x_reg_L0_22__retimed_I7645_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7645_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363;
	end
assign N13720 = x_reg_L0_22__retimed_I7645_QOUT;
reg x_reg_L0_22__retimed_I7642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7642_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383;
	end
assign N13712 = x_reg_L0_22__retimed_I7642_QOUT;
reg x_reg_L0_22__retimed_I7640_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7640_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307;
	end
assign N13706 = x_reg_L0_22__retimed_I7640_QOUT;
reg x_reg_L0_22__retimed_I7611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7611_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755;
	end
assign N13628 = x_reg_L0_22__retimed_I7611_QOUT;
reg x_reg_L0_22__retimed_I7610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7610_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339;
	end
assign N13626 = x_reg_L0_22__retimed_I7610_QOUT;
reg x_reg_L0_22__retimed_I7609_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7609_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242;
	end
assign N13624 = x_reg_L0_22__retimed_I7609_QOUT;
reg x_reg_L0_22__retimed_I7607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7607_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133;
	end
assign N13618 = x_reg_L0_22__retimed_I7607_QOUT;
reg x_reg_L0_22__retimed_I7606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7606_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851;
	end
assign N13616 = x_reg_L0_22__retimed_I7606_QOUT;
reg x_reg_L0_22__retimed_I7604_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7604_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173;
	end
assign N13610 = x_reg_L0_22__retimed_I7604_QOUT;
reg x_reg_L0_22__retimed_I7562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7562_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847;
	end
assign N13498 = x_reg_L0_22__retimed_I7562_QOUT;
reg x_reg_L0_22__retimed_I7561_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7561_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946;
	end
assign N13496 = x_reg_L0_22__retimed_I7561_QOUT;
reg x_reg_L0_22__retimed_I7560_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7560_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334;
	end
assign N13494 = x_reg_L0_22__retimed_I7560_QOUT;
reg x_reg_L0_22__retimed_I7554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7554_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222;
	end
assign N13478 = x_reg_L0_22__retimed_I7554_QOUT;
reg x_reg_L0_22__retimed_I7553_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7553_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322;
	end
assign N13476 = x_reg_L0_22__retimed_I7553_QOUT;
reg x_reg_L0_22__retimed_I7551_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7551_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088;
	end
assign N13470 = x_reg_L0_22__retimed_I7551_QOUT;
reg x_reg_L0_22__retimed_I7549_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7549_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357;
	end
assign N13465 = x_reg_L0_22__retimed_I7549_QOUT;
reg x_reg_L0_22__retimed_I7545_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7545_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478;
	end
assign N13455 = x_reg_L0_22__retimed_I7545_QOUT;
reg x_reg_L0_22__retimed_I7536_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7536_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479;
	end
assign N13432 = x_reg_L0_22__retimed_I7536_QOUT;
reg x_reg_L0_22__retimed_I7512_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7512_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940;
	end
assign N13366 = x_reg_L0_22__retimed_I7512_QOUT;
reg x_reg_L0_22__retimed_I7511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7511_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412;
	end
assign N13364 = x_reg_L0_22__retimed_I7511_QOUT;
reg x_reg_L0_22__retimed_I7494_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7494_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480;
	end
assign N13319 = x_reg_L0_22__retimed_I7494_QOUT;
reg x_reg_L1_15__retimed_I7474_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I7474_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735;
	end
assign N13263 = x_reg_L1_15__retimed_I7474_QOUT;
reg x_reg_L1_15__retimed_I7473_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I7473_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911;
	end
assign N13261 = x_reg_L1_15__retimed_I7473_QOUT;
reg x_reg_L1_22__retimed_I7470_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7470_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749;
	end
assign N13254 = x_reg_L1_22__retimed_I7470_QOUT;
reg x_reg_L0_22__retimed_I7467_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7467_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505;
	end
assign N13245 = x_reg_L0_22__retimed_I7467_QOUT;
reg x_reg_L0_22__retimed_I7466_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7466_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141;
	end
assign N13243 = x_reg_L0_22__retimed_I7466_QOUT;
reg x_reg_L0_22__retimed_I7465_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7465_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130;
	end
assign N13241 = x_reg_L0_22__retimed_I7465_QOUT;
reg x_reg_L0_22__retimed_I7463_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7463_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166;
	end
assign N13235 = x_reg_L0_22__retimed_I7463_QOUT;
reg x_reg_L0_22__retimed_I7458_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7458_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317;
	end
assign N13223 = x_reg_L0_22__retimed_I7458_QOUT;
reg x_reg_L0_22__retimed_I7455_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7455_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481;
	end
assign N13215 = x_reg_L0_22__retimed_I7455_QOUT;
reg x_reg_L0_22__retimed_I7434_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7434_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844;
	end
assign N13157 = x_reg_L0_22__retimed_I7434_QOUT;
reg x_reg_L0_22__retimed_I7433_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7433_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969;
	end
assign N13155 = x_reg_L0_22__retimed_I7433_QOUT;
reg x_reg_L0_22__retimed_I7432_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7432_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331;
	end
assign N13153 = x_reg_L0_22__retimed_I7432_QOUT;
reg x_reg_L0_22__retimed_I7429_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7429_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519;
	end
assign N13145 = x_reg_L0_22__retimed_I7429_QOUT;
reg x_reg_L0_22__retimed_I7423_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7423_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482;
	end
assign N13129 = x_reg_L0_22__retimed_I7423_QOUT;
reg x_reg_L0_22__retimed_I7402_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7402_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536;
	end
assign N13070 = x_reg_L0_22__retimed_I7402_QOUT;
reg x_reg_L0_22__retimed_I7401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7401_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277;
	end
assign N13068 = x_reg_L0_22__retimed_I7401_QOUT;
reg x_reg_L0_22__retimed_I7400_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7400_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155;
	end
assign N13066 = x_reg_L0_22__retimed_I7400_QOUT;
reg x_reg_L0_22__retimed_I7398_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7398_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236;
	end
assign N13060 = x_reg_L0_22__retimed_I7398_QOUT;
reg x_reg_L0_22__retimed_I7393_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7393_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345;
	end
assign N13048 = x_reg_L0_22__retimed_I7393_QOUT;
reg x_reg_L0_22__retimed_I7390_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7390_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483;
	end
assign N13040 = x_reg_L0_22__retimed_I7390_QOUT;
reg x_reg_L0_22__retimed_I7369_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7369_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983;
	end
assign N12979 = x_reg_L0_22__retimed_I7369_QOUT;
reg x_reg_L0_22__retimed_I7368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7368_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218;
	end
assign N12977 = x_reg_L0_22__retimed_I7368_QOUT;
reg x_reg_L0_22__retimed_I7367_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7367_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471;
	end
assign N12975 = x_reg_L0_22__retimed_I7367_QOUT;
reg x_reg_L0_22__retimed_I7364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7364_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794;
	end
assign N12967 = x_reg_L0_22__retimed_I7364_QOUT;
reg x_reg_L0_22__retimed_I7356_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7356_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484;
	end
assign N12945 = x_reg_L0_22__retimed_I7356_QOUT;
reg x_reg_L0_22__retimed_I7338_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7338_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734;
	end
assign N12895 = x_reg_L0_22__retimed_I7338_QOUT;
reg x_reg_L0_22__retimed_I7333_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7333_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485;
	end
assign N12881 = x_reg_L0_22__retimed_I7333_QOUT;
reg x_reg_L0_22__retimed_I7312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7312_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486;
	end
assign N12822 = x_reg_L0_22__retimed_I7312_QOUT;
reg x_reg_L0_22__retimed_I7298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7298_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575;
	end
assign N12781 = x_reg_L0_22__retimed_I7298_QOUT;
reg x_reg_L0_22__retimed_I7296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7296_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342;
	end
assign N12777 = x_reg_L0_22__retimed_I7296_QOUT;
reg x_reg_L0_22__retimed_I7293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7293_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150;
	end
assign N12769 = x_reg_L0_22__retimed_I7293_QOUT;
reg x_reg_L0_22__retimed_I7279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7279_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899;
	end
assign N12728 = x_reg_L0_22__retimed_I7279_QOUT;
reg x_reg_L0_22__retimed_I7278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245;
	end
assign N12726 = x_reg_L0_22__retimed_I7278_QOUT;
reg x_reg_L0_22__retimed_I7277_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7277_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390;
	end
assign N12724 = x_reg_L0_22__retimed_I7277_QOUT;
reg x_reg_L0_22__retimed_I7270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7270_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487;
	end
assign N12704 = x_reg_L0_22__retimed_I7270_QOUT;
reg x_reg_L0_22__retimed_I7256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7256_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488;
	end
assign N12663 = x_reg_L0_22__retimed_I7256_QOUT;
reg x_reg_L0_22__retimed_I7244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7244_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28];
	end
assign N12628 = x_reg_L0_22__retimed_I7244_QOUT;
reg x_reg_L0_22__retimed_I7242_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7242_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489;
	end
assign N12622 = x_reg_L0_22__retimed_I7242_QOUT;
reg x_reg_L0_22__retimed_I7231_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7231_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29];
	end
assign N12589 = x_reg_L0_22__retimed_I7231_QOUT;
reg x_reg_L0_22__retimed_I7230_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7230_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29];
	end
assign N12587 = x_reg_L0_22__retimed_I7230_QOUT;
reg x_reg_L0_22__retimed_I7228_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7228_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490;
	end
assign N12581 = x_reg_L0_22__retimed_I7228_QOUT;
reg x_reg_L0_22__retimed_I7216_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7216_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491;
	end
assign N12546 = x_reg_L0_22__retimed_I7216_QOUT;
reg x_reg_L0_22__retimed_I7205_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7205_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803;
	end
assign N12513 = x_reg_L0_22__retimed_I7205_QOUT;
reg x_reg_L0_22__retimed_I7204_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7204_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492;
	end
assign N12511 = x_reg_L0_22__retimed_I7204_QOUT;
reg x_reg_L0_22__retimed_I7183_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7183_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468;
	end
assign N12449 = x_reg_L0_22__retimed_I7183_QOUT;
reg x_reg_L0_22__retimed_I7181_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7181_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941;
	end
assign N12445 = x_reg_L0_22__retimed_I7181_QOUT;
reg x_reg_L0_22__retimed_I7173_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7173_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988;
	end
assign N12420 = x_reg_L0_22__retimed_I7173_QOUT;
reg x_reg_L0_22__retimed_I7172_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7172_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677;
	end
assign N12418 = x_reg_L0_22__retimed_I7172_QOUT;
reg x_reg_L0_22__retimed_I7171_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7171_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862;
	end
assign N12416 = x_reg_L0_22__retimed_I7171_QOUT;
reg x_reg_L0_22__retimed_I7153_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7153_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599;
	end
assign N12365 = x_reg_L0_22__retimed_I7153_QOUT;
reg x_reg_L1_22__retimed_I7147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7147_QOUT <= N12325;
	end
assign N12349 = x_reg_L1_22__retimed_I7147_QOUT;
reg x_reg_L1_22__retimed_I7141_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7141_QOUT <= N12309;
	end
assign N12333 = x_reg_L1_22__retimed_I7141_QOUT;
reg x_reg_L0_22__retimed_I7138_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7138_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452;
	end
assign N12325 = x_reg_L0_22__retimed_I7138_QOUT;
reg x_reg_L1_22__retimed_I7135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7135_QOUT <= N12295;
	end
assign N12317 = x_reg_L1_22__retimed_I7135_QOUT;
reg x_reg_L0_22__retimed_I7132_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7132_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781;
	end
assign N12309 = x_reg_L0_22__retimed_I7132_QOUT;
reg x_reg_L0_22__retimed_I7127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7127_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492;
	end
assign N12295 = x_reg_L0_22__retimed_I7127_QOUT;
reg x_reg_L1_22__retimed_I7126_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7126_QOUT <= N12274;
	end
assign N12291 = x_reg_L1_22__retimed_I7126_QOUT;
reg x_reg_L0_22__retimed_I7120_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7120_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985;
	end
assign N12274 = x_reg_L0_22__retimed_I7120_QOUT;
reg x_reg_L1_14__retimed_I7117_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I7117_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31];
	end
assign N12266 = x_reg_L1_14__retimed_I7117_QOUT;
reg x_reg_L1_16__retimed_I7114_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I7114_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006;
	end
assign N12259 = x_reg_L1_16__retimed_I7114_QOUT;
reg x_reg_L1_17__retimed_I7112_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I7112_QOUT <= N12076;
	end
assign N12254 = x_reg_L1_17__retimed_I7112_QOUT;
reg x_reg_L1_18__retimed_I7110_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I7110_QOUT <= N12071;
	end
assign N12249 = x_reg_L1_18__retimed_I7110_QOUT;
reg x_reg_L1_19__retimed_I7108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I7108_QOUT <= N12066;
	end
assign N12244 = x_reg_L1_19__retimed_I7108_QOUT;
reg x_reg_L1_20__retimed_I7106_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I7106_QOUT <= N12061;
	end
assign N12239 = x_reg_L1_20__retimed_I7106_QOUT;
reg x_reg_L1_21__retimed_I7104_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I7104_QOUT <= N12056;
	end
assign N12234 = x_reg_L1_21__retimed_I7104_QOUT;
reg x_reg_L1_22__retimed_I7102_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7102_QOUT <= N12051;
	end
assign N12229 = x_reg_L1_22__retimed_I7102_QOUT;
reg x_reg_L1_22__retimed_I7077_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7077_QOUT <= N11890;
	end
assign N12170 = x_reg_L1_22__retimed_I7077_QOUT;
reg x_reg_L1_22__retimed_I7076_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7076_QOUT <= N11888;
	end
assign N12168 = x_reg_L1_22__retimed_I7076_QOUT;
reg x_reg_L1_22__retimed_I7074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I7074_QOUT <= N11884;
	end
assign N12164 = x_reg_L1_22__retimed_I7074_QOUT;
reg x_reg_L0_17__retimed_I7039_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I7039_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654;
	end
assign N12076 = x_reg_L0_17__retimed_I7039_QOUT;
reg x_reg_L0_18__retimed_I7037_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I7037_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929;
	end
assign N12071 = x_reg_L0_18__retimed_I7037_QOUT;
reg x_reg_L0_19__retimed_I7035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I7035_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580;
	end
assign N12066 = x_reg_L0_19__retimed_I7035_QOUT;
reg x_reg_L0_20__retimed_I7033_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I7033_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983;
	end
assign N12061 = x_reg_L0_20__retimed_I7033_QOUT;
reg x_reg_L0_21__retimed_I7031_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I7031_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503;
	end
assign N12056 = x_reg_L0_21__retimed_I7031_QOUT;
reg x_reg_L0_22__retimed_I7029_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I7029_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772;
	end
assign N12051 = x_reg_L0_22__retimed_I7029_QOUT;
reg x_reg_L0_22__retimed_I6960_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6960_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29;
	end
assign N11890 = x_reg_L0_22__retimed_I6960_QOUT;
reg x_reg_L0_22__retimed_I6959_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6959_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67;
	end
assign N11888 = x_reg_L0_22__retimed_I6959_QOUT;
reg x_reg_L0_22__retimed_I6957_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I6957_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795;
	end
assign N11884 = x_reg_L0_22__retimed_I6957_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353 = !(a_exp[7] & a_exp[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355 = ((a_exp[4] & a_exp[3]) & a_exp[2]) & a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743 = !((a_exp[6] & a_exp[5]) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2355);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2353 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11743);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2376 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2395) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2384) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2404);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2389);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 = !(a_man[18] | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402 = !((((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381) | a_man[16]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2408) | a_man[15]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2393 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2402);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2387 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2378);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2523 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2514) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2526) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2518);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2516 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1] = !a_exp[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0] = !a_exp[0];
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[0]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2] = (!a_exp[2]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3] = !a_exp[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457 = !(a_exp[2] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2459);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5] = !a_exp[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[3] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2457);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451 = !(a_exp[4] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[5] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2451);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6] = (!a_exp[6]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7] = !a_exp[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444 = !(a_exp[6] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2449);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4] = (!a_exp[4]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2454;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[1]) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2464;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483 = !((((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2489) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[7] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2444);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2483 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2486) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__9) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__17);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N447));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448 = ((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[0] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N448;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11795 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__67;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427 = !a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 = !a_man[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 = !a_man[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 = !a_man[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 = !a_man[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 = !(a_man[16] & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3627 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 = !a_man[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 = !a_man[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3358 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3296 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3826 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 = !(a_man[17] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3668 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3282 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3504 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3829 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3416 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4007 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 = !(a_man[17] | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3457 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3283 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4023 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3626 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3458 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4011 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3849 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3629 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3214 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3809 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4022 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (a_man[19] & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054 = !(a_man[19] | a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3252 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4012 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3823 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3415 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841 = 1'B0 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N499;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7983} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7478};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7503 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[16]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3253 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3275 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3649 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3418 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3946 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3607 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3822 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3363 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3850 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3981 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3814 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3622 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3213 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 = !(a_man[17] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 = !((a_man[17] & a_man[16]) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3982 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3611 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3440 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3216 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3745 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3398 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3620 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4094 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3653 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3650 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3781 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3612 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3410 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3945 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783} = {1'B0, 1'B1} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N496};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N498;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7580 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N497) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7651;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] = !a_man[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3377 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3400 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3235 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3948 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3541 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4133 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3408 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3887 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3445 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3441 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3576 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3401 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3210 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3744 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3589 & a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 = !a_man[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4054);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3529 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4119 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16] = !(a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3606);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 = !a_man[13];
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6061} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6087};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6468} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6526};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N495} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[33]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7571};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7706} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7866} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7783};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7929 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3787 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4110 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4135 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3603 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3968 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3337 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3932 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3207 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3688 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3238 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3236 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3376 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4136 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3944 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3540 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637 = !a_man[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3563 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3323 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3915 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3848 | a_man[21]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3396 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3528 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6522} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6579};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888 = !a_man[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3361 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3919 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3750 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4049 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3710 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3928 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4092 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4122 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4132 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3322 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6116} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6200};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6549} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6482} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6070};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6257} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5773};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[32]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[32]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7988} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7645};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7599} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7460} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7886};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7654 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4125 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3929 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3902 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3935 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3767 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3864 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4063 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3729 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3939 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3480 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3970 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3560 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4109 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3936 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3742 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3336 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 = !a_man[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4093 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3715 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3845 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3508 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3725 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3987 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3743 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3885 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3920 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3930 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4048 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6576} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5825};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6143} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6173} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6326};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5740} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5768} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5798};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6291} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5840} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5807};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5995} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6448} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6371};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7862, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[31]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[31]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7677, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7468} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7725};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809} = {1'B0, N12416} + {1'B0, N12418} + {1'B0, N12420};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8006 = N12365 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3331 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3700 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3731 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3559 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3665 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3862 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3525 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3295 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3740 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3273 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3769 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4089 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3901 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3732 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N492 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3539 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4062 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747 = !a_man[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3886 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3512 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3342 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3646 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3300 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3523 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3788 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3872 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3984 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3686 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3716 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3727 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3844 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6170} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6310};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6198} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6225} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6252};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5792} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6137} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6165};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648 = !a_man[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5765} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5795};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[13];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5744} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6465};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6514} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6546} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6028};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[29]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6214} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6182} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5731};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7941, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7803} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[30]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[30]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572} = {1'B0, N12511} + {1'B0, N12513};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022} = {1'B0, N12445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7892} + {1'B0, N12449};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3516 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3497 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3531 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3359 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3455 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3663 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3320 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3537 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4002 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3566 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3883 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3699 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3532 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N491 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3334 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3861 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 = !a_man[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3479 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4031 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3868 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3561 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3232 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3828 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4040 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3381 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3462 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3579 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3270 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3306 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3318 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3436 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6223} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6421};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[12];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6187} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5877} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5907};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3687 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3305 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4070 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3768 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3437 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4027 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3316 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3582 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[18] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3673 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3783 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3478 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3513 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3524 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3645 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5934} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5823} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5850};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6119} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6496} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5980};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6278} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6308};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 = !a_man[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3271 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3834 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3395 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3669 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3360 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3965 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3628 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430 = !(a_man[19] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3430 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4115 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3258 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3380 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4000 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4033 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4043 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3231 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6041};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6247} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6338} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6366};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6418} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6561} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6074};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6245} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6358} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6010} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5869};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[29], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[28]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6056} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6405} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6434};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888} = {1'B0, N12587} + {1'B0, N12589};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674} = {1'B0, N12546} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7888};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8018} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7572};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3288 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3324 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3237 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4088 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3249 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3454 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4045 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3255 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3330 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3805 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3705 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3365 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3684 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3496 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3325 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N490 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4061 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3662 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[11];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5848} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5875} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5904};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6397} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5999} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5762};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6390, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5932} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6307} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6453};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[10];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698 = !a_man[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4055 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4001 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3633 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3755 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3459 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4090 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3764 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3417 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3827);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3956 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3908 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3244 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3988 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4113 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3803 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3835 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3841 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3964 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6276} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6534};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5937} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6017} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5933};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5961} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5989} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6058};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5777} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6140} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6375} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6517};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5899, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6575} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5965} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5822} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6197};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]} = {1'B0, N12724} + {1'B0, N12726} + {1'B0, N12728};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965} = {1'B0, N12628} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[28]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776} = {1'B0, N12581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7965};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7700} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7674};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3657 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4018 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4050 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3882 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3979 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3247 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3842 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4078 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4057 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3599 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4095 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3476 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3287 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4051 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N489 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3859 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3453 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[9];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6504} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6419} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6449};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6409, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6218} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6203} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5951} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6329};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11689;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6304} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6335} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6363};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 = !a_man[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 = !a_man[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3598 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3219 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3983 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3685 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3355 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3947 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3549 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3502 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4041 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3672 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3584 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3704 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3391 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3425 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3433 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3555 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6333} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5780};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[8];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6071} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5908} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6127};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3911 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3397 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3804 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3423 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3907 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4076 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3254 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3884 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3556 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3215 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3830 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3756 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3706 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3790 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3906 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3597 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3634 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3640 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3763 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5873} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6153};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6109} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6477} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6394};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6003} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6123} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6500};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5900} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5930} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5958};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6097} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5987} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6014};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5746} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6489} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6380};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5827} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6436};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5919, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5734} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6581} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6089} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5842};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530} = {1'B0, N15285} + {1'B0, N15287} + {1'B0, N15289};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6342, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6150} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5885} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6261} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6030};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]} = {1'B0, N12777} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5854} + {1'B0, N12781};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[27]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[27]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876} = {1'B0, N12622} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7420};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7917} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7776};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3819 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3846 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3362 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3683 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3778 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3978 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3642 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3855 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3392 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3754 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3535 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3690 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3267 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4017 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3847 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N488 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3661 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3246 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6361} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6392} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6416};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6039} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5923} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6283};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6558} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6445} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6475};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 = !a_man[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 = !a_man[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 = !a_man[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6389};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5929} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6098};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6194} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6531} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5728};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5800} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6297};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6471, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6277} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5890} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6013} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6266};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[7];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5749} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6501} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5725};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6551} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6190} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5814};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5983, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5794} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6393} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5782} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5903};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105} = {1'B0, N12975} + {1'B0, N12977} + {1'B0, N12979};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]} = {1'B0, N12769} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6294} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6530};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[26]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[26]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982} = {1'B0, N12663} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7508};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7634} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7511} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7876};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3326);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3402 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 = a_man[22] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3467;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2681} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2704};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748, N15860} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2772} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2711};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2784} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2748} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2638};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2816} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2804} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2879};
assign {N15894, N15886} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2746} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2694};
assign {N15865, N15853} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2630} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2642} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2870};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889, N15878} = {1'B0, N15894} + {1'B0, N15860} + {1'B0, N15865};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2670} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2768};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2659} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2829};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2593} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2624};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2713} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2699};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2701} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2776} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2812};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11653;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2666} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2785} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2635};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2679} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2782} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2736};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2798} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2644} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2614};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2712} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2780} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2602};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2845} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2655};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2854} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2671} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2844};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2825} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2839};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2885) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2790;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880, N15996} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2611} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2708};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2587} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2880};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2787} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2754} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2604};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2709} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2691};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2742} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2647};
assign {N16030, N16016} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2851} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2820} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2806};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695, N16042} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2859} + {1'B0, N16030} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2665};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2865} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2695} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2683};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2673} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2834} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2830};
assign {N16022, N16008} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2619} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2650} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2794};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841, N16034} = {1'B0, N15996} + {1'B0, N16022} + {1'B0, N16042};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2637);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2788} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2878};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2888);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2609} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2595};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702, N16079} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2685} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2680};
assign {N16014, N16003} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2702};
assign {N16115, N16101} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2715} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2732};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846, N16128} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2856} + {1'B0, N16115} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2819};
assign {N16020, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2872} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2846} + {1'B0, N16003};
assign {N16107, N16095} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2862} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2868} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2684};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660, N16120} = {1'B0, N16107} + {1'B0, N16079} + {1'B0, N16128};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2747);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2698 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2648);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2779};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2616} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2636};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11697);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2631 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2629} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2822};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2763} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2626};
assign {N16087, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2590} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2770} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2656};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11662} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2675};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11670);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2764) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2895)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2815) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2739));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2628 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2586) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2814 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2882)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2723) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2869)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2697) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2842));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2589 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2800);
assign {N16099, N16089} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2727} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2721};
assign {N16126, N16113} = {1'B0, N16101} + {1'B0, N16099} + {1'B0, N16095};
assign N16085 = !N16126;
assign N16121 = !((N16120 & N16085) | ((!N16120) & N16126));
assign {N16105, N16093} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2726} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2615} + {1'B0, N16089};
assign N16116 = !N16105;
assign N16123 = !(N16116 & N16113);
assign N16084 = !(N16116 | N16113);
assign N16075 = !N16084;
assign N16111 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2745 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2863) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2797);
assign N16082 = !((N16087 & N16093) | N16111);
assign N16108 = !(N16087 | N16093);
assign N16091 = !(N16108 | N16082);
assign N16080 = !(N16105 | N16113);
assign N16119 = !((N16075 & N16123) | N16091);
assign N16104 = !(N16080 | N16119);
assign N16102 = N16126 | N16120;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576 = ((!N16121) & (!N16104)) | (!N16102);
assign {N16039, N16027} = {1'B0, N16014} + {1'B0, N16016} + {1'B0, N16008};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652 = N16039 ^ N16034;
assign N16005 = !N16020;
assign N16010 = !(N16005 & N16027);
assign N16029 = !(N16005 | N16027);
assign N16017 = !N16029;
assign N16032 = N16020 ^ N16027;
assign N15993 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2837;
assign N16001 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2689 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2576);
assign N16012 = !(N15993 & N16001);
assign N16025 = !(N16020 | N16027);
assign N16040 = !((N16017 & N16010) | (N15993 & N16001));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871 = (N16012 & N16032) | N16025;
assign N15997 = !(N16039 | N16034);
assign N16038 = !N15997;
assign N16019 = ((!N16040) & (!N16025)) | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749 = !(N16038 & N16019);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2841 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2832);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2720;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2896 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2741);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2861;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2817 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2658);
assign {N15858, N15845} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2894} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2632} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2774};
assign {N15883, N15873} = {1'B0, N15886} + {1'B0, N15858} + {1'B0, N15853};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852 = N15883 ^ N15878;
assign {N15863, N15851} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2802} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2591} + {1'B0, N15845};
assign N15861 = !N15863;
assign N15867 = !(N15861 & N15873);
assign N15885 = !(N15861 | N15873);
assign N15875 = !N15885;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710 = N15863 ^ N15873;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729 ^ N15851;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2678;
assign N15856 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2729 | N15851);
assign N15888 = !N15856;
assign N15870 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893) | N15856;
assign N15854 = !N15873;
assign N15881 = !(N15863 | N15873);
assign N15871 = !((N15875 & N15867) | (N15888 & N15870));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 = (N15861 & N15854) | N15871;
assign N15849 = !(N15883 | N15878);
assign N15869 = !N15849;
assign N15848 = ((!N15871) & (!N15881)) | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703 = !(N15869 & N15848);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2889 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2778);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign N15963 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777);
assign N15934 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777;
assign N15944 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809, N15952} = {1'B0, N15934} + {1'B0, N15963} + {1'B0, N15944};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809);
assign N15832 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2696;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2668 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2809;
assign {N15947, N15939} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2831} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2853} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2706};
assign N15929 = !N15952;
assign N15933 = !(N15929 & N15947);
assign N15959 = !N15947;
assign N15940 = !(N15952 & N15959);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625 = N15952 ^ N15947;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813 = N15939 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2599;
assign N15942 = !(N15939 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2849);
assign N15949 = !N15942;
assign N15935 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813) | N15942;
assign N15957 = !(N15952 | N15947);
assign N15936 = !((N15940 & N15933) | (N15949 & N15935));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2811 = (N15929 & N15959) | N15936;
assign N15834 = ((!N15936) & (!N15957)) | (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2769);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2803 = !(N15832 & N15834);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2588 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2848));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24] = (!N15271) ^ N14301;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[24];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24] = !(N13060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3674 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3343 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3406 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3438 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3225 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3266 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3374 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3572 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3228 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3728 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3449 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3926 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3274 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3800 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3616 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3439 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N486 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3245 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3776 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3866 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3573 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3798 | a_man[20]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3261 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3592 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N457;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154 = !(N13235 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23] = N14406 ^ N14408;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219 = !(N13060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341 = !(N13235 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[22] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2634) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2625;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367 = !N14435;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072 = !(N13060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3753 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3711 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3310 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3918 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3373 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917 = !(a_man[21] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3991 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3917 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N456;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274 = !(N13470 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5072} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5274};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5219} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5349};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010} = {1'B0, N12822} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[24]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 = !(a_man[18] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3617 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3647 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3475 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3574 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3777 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3434 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3931 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3581 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3656 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4129 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3874 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3548 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3481 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3997 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3818 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3648 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N487 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3451 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3977 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6012} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6124} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6183};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3995);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4128 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3951 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3782 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3477 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4085 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3746 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3429 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3489 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3348 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3292 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3383 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3500 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4127 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3220 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3226 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3354 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6264} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5956} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5985};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6151} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6038} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6067};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6568} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6461};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[6];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6209} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6235} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6093};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6095} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5973} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6474};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6155, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5969} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6063} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6565} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6439};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5747} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6528};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5808} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5835} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6555};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5879} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6253};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 = !(a_man[16] & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3293 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3720 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3545 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3485 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3379 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3998 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3680 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3338 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3394 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3638 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3315 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3873 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3409 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3810 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3957 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3909 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4020 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3719 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3749 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3758 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3878 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5982} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6378} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5922};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5726} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6493} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5778};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6367} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5894} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6269};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6331, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6141} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5863} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5874} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6236};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4025 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3999 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3925 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3748 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4098 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3578 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3268 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3879 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3542 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3522);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4077 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3621 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4008 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4116 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3291 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3924 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3952 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3959 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4084 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5888} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6414} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5914};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6009} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6034} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6065};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[5];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6321} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6180} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6232};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6387} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6286} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5896};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[4];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6092} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6121};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6206} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6262} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6290};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6442} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6473} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5860};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5790} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6272} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5803};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5786} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5769} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6145};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6479} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6005} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5990};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5986} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6350} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6364};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5844, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6519} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5751} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5766};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857} = {1'B0, N13153} + {1'B0, N13155} + {1'B0, N13157};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6536, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6345} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6078} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5954} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6456};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169} = {1'B0, N13066} + {1'B0, N13068} + {1'B0, N13070};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]} = {1'B0, N12967} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6043} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6169};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]} = {1'B0, N12895} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6360} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6105};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[24]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[24]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459} = {1'B0, N12704} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7530} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7795};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[25]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[25]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7719} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7722} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7982};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4099 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3596 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3519 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3340 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3277 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3941 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4112 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3801 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3472 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4064 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3551 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3675 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3208 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3608 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3757 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3891 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3789 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3707 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3821 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3518 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3546 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3552 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3679 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6035);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6438} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6002} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6469};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6407} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6148} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6303};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6334} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6554} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6163} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6066};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6130, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5940} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6160} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6523} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6539};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[3];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5972} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5804} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5858};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6494} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6525} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5916};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5775} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6553} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5831};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5917} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5809} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6292};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5944} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5886} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5745};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6196} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6184} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6572};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5847} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6179} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6545} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6053};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6505, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6317} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6048} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6033} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6427};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031} = {1'B0, N13241} + {1'B0, N13243} + {1'B0, N13245};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]} = {1'B0, N13048} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5857};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[23]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8010} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7659} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7874};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7585} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7937} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7459};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4056 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3806 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3269 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3206 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3233 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3272 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3996 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4106 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3372 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3961 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3949 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3990 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3241 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3721 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3466 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4004 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3594 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3405 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3234 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N485 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3975 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3571 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195 = !(N13235 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2601) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2813;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260 = !(N13060 | N15245);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127 = !(N13470 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5195} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5127};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318 = !(N13470 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387 = !(N13235 | N15245);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2703 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2667;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115 = !(N13060 | N15230);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5387} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5318} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5115};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3547 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3577 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3666 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3250 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3452 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3738 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4035 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3713 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4105 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4071);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3796 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3510 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N455;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401 = !(N13465 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5401} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5332} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5171};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5244} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5272} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5392};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471} = {1'B0, N12881} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[23]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[23]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3276 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3312 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4068 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4006 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3905 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3595 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3265 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3863 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3736 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3464 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3942 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3693 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3486 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3583 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3503 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3619 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3311 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3341 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3349 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3471 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6446);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6062} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6488} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6088};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5724} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6215} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6309};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6242} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6463} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6084} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6559};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6412, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6222} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6444} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6430} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5957};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[2];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6459} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6146} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6318};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6229} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6406};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6118} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6287};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6577} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5824};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6346} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6205};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6086} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5732} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6483};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5946, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5755} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6072} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5978} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6450};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738} = {1'B0, N13494} + {1'B0, N13496} + {1'B0, N13498};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833} = {1'B0, N13364} + {1'B0, N13366} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5927};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]} = {1'B0, N13145} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6019} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6031};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3601 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3938 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3966 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3799 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3898 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4104 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3760 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3793 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3501 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3972 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3520 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3807 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3388 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3205 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3967 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N484 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3775 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3371 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552} = {1'B0, N12945} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[22]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[22]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7471} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7686};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7606} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7533} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7565};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4079 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3726 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3345 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3378 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4091 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3536 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3837 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3511 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3897 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3297 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3737 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904 = !(a_man[20] | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3538);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3870 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3904 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3588 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3303 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N454;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185 = !(N13745 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249 = !(N13465 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5173 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2627 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2852;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5305 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237 = !(N13235 | N15230);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196} = {1'B0, N15281} + {1'B0, N13610} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5237};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5249} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5268};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379 = !(N13745 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106 = !(N13465 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4072 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4111 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3488;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3209 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3329 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3635 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3304 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3696 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3610 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4024 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3854 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4015 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3333 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3655 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3670 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3702 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3385 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4029 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N453;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310 = !(N13925 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5106} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5310};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5254} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5066};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5143} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5317} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5288};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[22]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[22]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3413 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3985 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4126 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4038 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3867 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3605 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3332 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3703 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3389 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3994 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3664 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3808 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3301 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3639 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3259 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3741 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4134 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[17] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3382 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3294 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3407 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4037 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4069 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0] = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4081 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3264 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[33] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5992);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5830} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5856} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6000};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6177} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5843} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6487};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5774} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6102} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5996} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6467};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6322, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6133} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5962} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5866};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6580} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5968} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5883};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6052} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5743} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5915};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5736} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6120};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[1];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6403);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6172} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6201};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6126};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6027} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5941} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5802};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6001} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6377} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6498};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6339, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6147} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5981} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6372} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6359};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511} = {1'B0, N13624} + {1'B0, N13626} + {1'B0, N13628};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112} = {1'B0, N13476} + {1'B0, N13478} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5836};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]} = {1'B0, N13223} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6299} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5833};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (a_man[16] & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3352 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3860 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3735 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3765 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3444 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3448 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4032 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3593 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3697 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3895 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3553 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4044 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3586 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3772 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3313 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3347 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[16]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3869 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3463 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3364 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3602 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4124 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3937 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3766 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N483 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3569 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4103 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627} = {1'B0, N13040} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[21]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7767} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7817} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7552};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7957} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7744} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7663};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6547} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6391} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6011} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5901};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5851, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6527} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5882} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5870} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6258};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[0];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2777 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6227} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6567} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6256};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6425} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6515} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6344};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6502} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5905} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6296};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6316} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6373};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6108) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6550;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6486} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6401};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6518} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6016} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6396};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6246, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6057} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5887} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6263} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6275};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037} = {1'B0, N13780} + {1'B0, N13782} + {1'B0, N13784};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023} = {1'B0, N13616} + {1'B0, N13618} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6226};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5738} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6112};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3309 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4108 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4074 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3419 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3534 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3557 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4075 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493 = !((a_man[18] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[16] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3387 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3493 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3695 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3350 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3482 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4021 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3567 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4039 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3794 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[17]);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3689 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3393 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3922 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3734 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3558 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N482 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3370 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3894 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709} = {1'B0, N13129} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[20]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2580 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2893;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2690 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2710;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5383, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5307} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5281} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5347} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5214};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3526 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3432 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3871 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3903 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3943 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3426 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4030 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3492 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3570 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3795 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3279 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3824 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3568 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3229 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3614 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4059 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3447 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3460 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3499 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4118 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3832 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N452;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094 = !(N15238 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355 = !(N13925 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081 = !(N13745 | N15245);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5150 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5081} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5355} + {1'B0, N13917};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5094} + {1'B0, N13712} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5189};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5089 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5159 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5297 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326} = {1'B0, N13751} + {1'B0, N13753} + {1'B0, N13755};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3671 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3701 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3390 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4120 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3654 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3221 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3833 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3284 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3840 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3811 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3792 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3623 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3367 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3876 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (a_man[17] & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4058 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3858 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3240 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3256 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3290 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3914 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3631 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N451;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220 = !(N14060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5217, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5145} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5068} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5339};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286 = !(N15238 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263} = {1'B0, N13889} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5220} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5286};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5363 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231 = !(N13745 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164 = !(N13925 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5231} + {1'B0, N13720} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5164};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5337} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5326} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5137};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5343} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5358} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5167};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5400} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5208} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5196};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5228} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5376} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5213};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[21]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[21]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7838} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7627} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7902};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7961} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7770};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5920} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6410} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5812};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5760, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6435} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5793} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5779} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6167};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6024} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6162};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2705 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6543} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5924} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5938};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6079} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6049} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5997};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5881} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5912} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5966};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5947);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6106} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5799} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5939};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5816} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6192} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6298};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6152, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5967} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6280} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6188} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5797};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5826} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6138} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5853};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6566} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5829} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6204};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6532, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6343} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6563} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6171} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6075};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950} = {1'B0, N13944} + {1'B0, N13946} + {1'B0, N13948};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415} = {1'B0, N13759} + {1'B0, N13761} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6139};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6511} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5741} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6023};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4080 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3431 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3328 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3356 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3260 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3636 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3771 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4123 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3285 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3491 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4082 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3752 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3976 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3761 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3442 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3366 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3839 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3708 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3587 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3543 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3969 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4130 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3718 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3533 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3357 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N481 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4100 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3694 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787} = {1'B0, N13215} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[19]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270 = !(N13745 | N15230);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141 = !(N15238 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073 = !(N14060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5141} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5270} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5073};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2603 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2752;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5200 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5135 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5206 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291} = {1'B0, N14079} + {1'B0, N14081} + {1'B0, N14083};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5364} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5175} + {1'B0, N13706};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5398 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262 = !(N14060 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4067 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3785 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4042 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3461 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3498 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4026 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3550 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3446 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3953 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3632 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4013 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3414 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4101 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3494 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3412 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4097 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3351 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3658 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3971 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3986 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4019 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3709 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3421 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N450;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197 = !(N14214 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[23]);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5262} + {1'B0, N14024} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5197};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5124 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2766 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2610;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5391 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5330 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123} = {1'B0, N14071} + {1'B0, N14073} + {1'B0, N14075};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5198} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5345} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5291};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2749 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2795;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5225, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5152} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5242} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5314} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5177};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3724 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3992 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3319 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3257 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3289 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3857 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3893 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3384 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4117 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3239 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3751 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3422 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3815 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3530 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3506 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3212 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3211 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3889 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3989);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3923 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3243 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3770 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3786 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3820 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3507 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3218 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 = !float_div_cynw_cm_float_rcp_E8_M23_3_inst_N449;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129 = !(N14209 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5372, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5298} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5384} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5110} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5247};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5129} + {1'B0, N13867} + {1'B0, N13869};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342 = !(N14214 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5176);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5389, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5313} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5191} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5256} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5325};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5342} + {1'B0, N13883} + {1'B0, N13885};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5157} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5099} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5246};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5128} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5075} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5275};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5118} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5321} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5263};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5149} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5283} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5295};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5090} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5104} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5239};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5155} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5312} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5299};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[19]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[19]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7924} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7709} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7575};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[20]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[20]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7497} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7557} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7868};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11728 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6484} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5759};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6564} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6369} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6400};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6096} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5737} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6476};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6315} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5723} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6080};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6540} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6455} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6311};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6341} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6512} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6424};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5988} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6365} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6490};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5872} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6091} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6458} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6472};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6040, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5855} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6548} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6454} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6060};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327} = {1'B0, N13767} + {1'B0, N13769} + {1'B0, N13771};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6037} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6516} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6415};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3424 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3784 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3399 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3404 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4053 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4086 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3625 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3317 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3618 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3921 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4014 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3281 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3875 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3227 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3660 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3912 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3739 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4096 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3637 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4137 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3856 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3344 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3585 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3562 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3927 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3515 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3327 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4087 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N480 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3892 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3490 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864} = {1'B0, N13319} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[18]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8001} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7787} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7434};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7980} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7771} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7969};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6356);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11719 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6076} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6219};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6282} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5789};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5784} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6111} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6004} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5876};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6437, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6248} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5970} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5984} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6362};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230} = {1'B0, N13931} + {1'B0, N13933} + {1'B0, N13935};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5950} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6420} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6327};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3565 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3580 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3248 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3853 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3880 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3450 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3958 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3933 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3717 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3816 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4010 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3677 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3960 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3590 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3779 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3428 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3505 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3242 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4003 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3722 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3308 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4052 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3881 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N479 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3692 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3280 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945} = {1'B0, N13432} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[17]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388 = !(N14214 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5116 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181 = !(N15238 | N15230);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107} = {1'B0, N14030} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5388} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5181};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320 = !(N14209 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11739);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2871 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2652;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5236 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5397, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5322} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5096} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5233};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5205, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5132} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5368} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5101} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5301};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250} = {1'B0, N14014} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5320} + {1'B0, N14018};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5179} + {1'B0, N13859} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5328};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5166 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5380, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5304} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5222} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5360};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5306 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174 = !(N14209 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5367);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086} = {1'B0, N14166} + {1'B0, N14168} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5174};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5374 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5168 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5238 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278} = {1'B0, N14202} + {1'B0, N14204} + {1'B0, N14206};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5354} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5163} + {1'B0, N14002};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5123} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5269} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5139};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5395} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5303} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5113};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5223} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5083} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5370};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[18]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[18]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7457} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7864} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7520};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7649} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7984} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7450};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3564 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4065 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3899 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3652 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3681 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3723 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3791 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3838 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3940 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3469 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3514 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3613 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3813 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3468 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3974 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3298 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3643 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3691 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3224 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3517 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3222 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4046 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3973 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3910 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3802 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3521 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4034 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3852 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3682 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N478 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3487 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4009 & a_man[22]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11661 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5935} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6103} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6022};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6158} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5964} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5994};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5911} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6542} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6161};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6134} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6047} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6191};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6051} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5801} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6284};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6347, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6156} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6382} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5767};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11708 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6538} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5815};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5897);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5906} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5849} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6462};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5756} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6422} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6452};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6305);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6398} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6562} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6481};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5733} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6509} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5787};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5739} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6224} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6115};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6176} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6428} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5943};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5859, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6537} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5891} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6267} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6142};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764} = {1'B0, N14087} + {1'B0, N14089} + {1'B0, N14091};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]} = {1'B0, N13727} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5952} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6230};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890 = N13455 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5169, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5093} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5344} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5147};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5091 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071} = {1'B0, N14316} + {1'B0, N14318} + {1'B0, N14320};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386} = {1'B0, N14006} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5146} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5278};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5120} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5250} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5402};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5088 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5186, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5114} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5156} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5226} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5085};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5160 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5293 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5365 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5294);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259} = {1'B0, N14284} + {1'B0, N14286} + {1'B0, N14288};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234} = {1'B0, N14158} + {1'B0, N14160} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5334};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209} = {1'B0, N13849} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5107} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5309};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5080} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5285} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5230};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5092} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5378} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5184};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[16]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7890} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7945} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7806};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5203} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5257} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5351};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[17]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[17]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7578} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7561};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757 = (!N13455) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 = !((a_man[17] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3346 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3676 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3299 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3733 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3443 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3473 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3369 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3223 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3759 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3913 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3307 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3403 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3609 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3262 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3335 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4073 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3825 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4102 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3483 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3955 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773 = !((a_man[16] & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3641) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4036 & a_man[18]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3624 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3773 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2381 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3714) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3600 & a_man[19]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3314 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3411) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3836 & a_man[20]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3651 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3474 & a_man[21]));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N477 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3278 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3427) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3812 & a_man[22]));
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6352} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5976} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5864};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6521, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6332} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6552} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6064} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6320};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046} = {1'B0, N14230} + {1'B0, N14232} + {1'B0, N14234};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6233} + {1'B0, N13907} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5764};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487} = {1'B0, N13735} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7618} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7757} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[16]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7597} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7655};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5282 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5078 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5216 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5221);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390} = {1'B0, N14402} + {1'B0, N14398} + {1'B0, N14400};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5315, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5240} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5276} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5348} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5210};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218} = {1'B0, N14174} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5125} + {1'B0, N14178};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5086} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5292} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5234};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5209} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5359};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7487} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[15]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8005} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7675} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7763};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11706 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6132} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6270};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5852);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6216} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6018} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6042};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6524} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5806};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6189} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6157} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6073};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6181} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6413} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6036};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6508} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6492} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6239} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6007};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6032, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5846} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6441} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5834} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5955};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]} = {1'B0, N14038} + {1'B0, N14040} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6046};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5357 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5108, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5373} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5131} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5267};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5252, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5180} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5403} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5136} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5335};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199} = {1'B0, N14324} + {1'B0, N14326} + {1'B0, N14328};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5271} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5259} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5071};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5386} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5192};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[14]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[15]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7601} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7861};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11693 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5730} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5867};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6100} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6243} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6244};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6260);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5813} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5754} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6503};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5785} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6535} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6560};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6101} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5758} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6136};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6195} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6557} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5928} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6069};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6208, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6021} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5753} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6386} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6131};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]} = {1'B0, N14182} + {1'B0, N14184} + {1'B0, N14186};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5069 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5148);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5201 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5280 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5194, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5251} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5393};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329} = {1'B0, N14419} + {1'B0, N14421} + {1'B0, N14423};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346} = {1'B0, N14278} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5064} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5390};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5082} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5218} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5366};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[13]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[14]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7811} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7964};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6186} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6328};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11688 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5841} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6574} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6055};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6255} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5993} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6480} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6513};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5895, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6571} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6302} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6447} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5818};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]} = {1'B0, N14292} + {1'B0, N14294} + {1'B0, N14296};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5074);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5340, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5266} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5187} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5258} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5122};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140} = {1'B0, N14382} + {1'B0, N14384} + {1'B0, N14386};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5211} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5199} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5346};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[12]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[13]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8024} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7442};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6240} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6154} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6295};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5810);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6268} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6213} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6128};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5839} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6085} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6464} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6433};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5960, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5772} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6370} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6026} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5880};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]} = {1'B0, N14390} + {1'B0, N14392} + {1'B0, N14394};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5865} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5811} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5838};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2773 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5781} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5921};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6417} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5931} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6388};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6404, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6212} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5948} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5979} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6324};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]} = {1'B0, N14469} + {1'B0, N14471} + {1'B0, N14473};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5235, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5311} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5112} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5243};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5207 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5381} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5178};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5336);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5153, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5077} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5327} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5087} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5121};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]} = {1'B0, N14374} + {1'B0, N14376} + {1'B0, N14378};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[10]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]} = {1'B0, N14260} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5329} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5140};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[11]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[11]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7832} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7648};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7622} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[12]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7550};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6217);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5761);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11669 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6234} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6383};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5750} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5892} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5776};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6357, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5898} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6306} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6273};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]} = {1'B0, N14505} + {1'B0, N14507} + {1'B0, N14509};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5134 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5261);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5165} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5302};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5399 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5188);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5289} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5158};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5097} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5369} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5323};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[9], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[8]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5133} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5356} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5279};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[9]} + {1'B0, N14370};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[10]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7429} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7753};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6325} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6265} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6293};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6149} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6228} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5742};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[8], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[7]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5821} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5791} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6164};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960} = {1'B0, N14454} + {1'B0, N14456} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[8]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7643} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[9]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7851};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5918} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5949};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6353} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6374} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6451};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[7], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[6]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6529} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6117} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6495};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437} = {1'B0, N14487} + {1'B0, N14489} + {1'B0, N14491};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995} = {1'B0, N14339} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7857} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7960};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N11660 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5889} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5861} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5977};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[5]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5884} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5963} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6340};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7451, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7542} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[6]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[6]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592} = {1'B0, N14441} + {1'B0, N14443} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7437};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5117);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6379} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6408};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N2876 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6578);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6122);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5975 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5971} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6029};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6349} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6432} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6104};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5], float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6485} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6185} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5998};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5324 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7667, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7640} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[5]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[5]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802} = {1'B0, N14479} + {1'B0, N14481} + {1'B0, N14483};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5248 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N5382);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7884, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[4]};
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016} = {1'B0, N14515} + {1'B0, N14517} + {1'B0, N14519};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802;
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7748, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[4]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7745};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444 = !(N14494 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[3]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[3]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533);
assign {float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562, float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417} = {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[2]} + {1'B0, float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[2]};
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909 = !(((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6570 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6301) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6533) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N6077);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7909 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7417);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7562 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7823);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7998 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7532) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8012);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7605 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7797) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7837)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7963) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7612));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936 = !(N14494 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8016);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989 = !((N14465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7444) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7936);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7721) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7989)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7535) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7802));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7939 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7592);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7670 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7991) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7849);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7635) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7973)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7724) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7995));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7514 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7780);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7583 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7916) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7777);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7564) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7800)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7919) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7570));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7703 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7971);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7948 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7826) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7699);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540 = ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7486) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7474)) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7491) & (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7761));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7895 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7545);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419 = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7754 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7540) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7615;
assign N14535 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7419 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7824) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7679 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7952)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558 = !N14535;
assign N14543 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7558 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7481) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7464 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7733)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747 = !N14543;
assign N14551 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7747 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7750) | (!(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7869 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7524)));
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590 = !N14551;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7653 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7927;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7488) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7439 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7712;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7807) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7501 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7844;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7521) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7906 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7631;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7840) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7415 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7690;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7553) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7476 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7821;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7875) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7880 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7610;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7586) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7664 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8013;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7914) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7447 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7799;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7614) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7853 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7589;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7942) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7638 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7992;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7646) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7425 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7778;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7976) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7829 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7568;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7683) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7620 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7968;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8009) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8022 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7758;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7716) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7809 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7543;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7736 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7418) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7735 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7911);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7749 = N12365 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7947;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7452 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8003 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7732;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7781 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7789 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7523;
assign N16185 = !(N15293 & N12259);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831 = (!N13254) | (N15293 & N12259);
assign N16186 = !N12254;
assign N16199 = !((N16185 & N13254) | N16186);
assign N16197 = !N12349;
assign N16203 = !(N16197 | N16199);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588 = (!N12349) | (N12254 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831);
assign N16201 = !N12249;
assign N16190 = !(N16201 | N16203);
assign N16194 = !N12333;
assign N16193 = !(N16194 | N16190);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608 = !N16193;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7492 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7926 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7582;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899 = (!N12317) | (N12244 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608);
assign N16169 = !N12234;
assign N16171 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899 | (!N12239));
assign N16168 = !(N16169 | N16171);
assign N16165 = !(N12291 | N16168);
assign N16167 = !N12229;
assign N16173 = !(N16167 | N16165);
assign N16162 = !((N12229 | N12291) | N16168);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834 = !N16171;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39] = !(N16162 | N16173);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7985 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7769 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7499);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896 = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_N4114 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3954);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N3896 | a_man[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N500 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7629;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7772 = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7894) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7904;
assign x[22] = (N12170 & N12164) | (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[39] & N12168);
assign N14526 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7834 ^ N12234;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38] = !N14526;
assign x[21] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[38]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7899) ^ N12239;
assign x[20] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[37]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7608) ^ N12244;
assign x[19] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[36]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7588) ^ N12249;
assign x[18] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[35]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7831) ^ N12254;
assign x[17] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[34]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33] = (!N15293) ^ N12259;
assign x[16] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[33]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32] = (!N13261) ^ N13263;
assign x[15] = (N12168 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[32]) | ((!N12168) & N12170);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[31] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7728) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7465;
assign x[14] = (N12168 & N12266) | ((!N12168) & N12170);
assign N14556 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7820 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7813;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30] = !N14556;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[13] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[30]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7567) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7546;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[29]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7579) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7896;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[28]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7856) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7623;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[27]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7794) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7972;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[26]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7996) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7704;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[25]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7847) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7430;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[24]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7979) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7782;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[23]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7756) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7515;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[22]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7798) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7858;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[21]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7500) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7593;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[20]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7462) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7940;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[19]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18] = (!float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7702) ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7668;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[18]) | ((!N11888) & N11890);
assign N14562 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_N7590 ^ float_div_cynw_cm_float_rcp_E8_M23_3_inst_N8017;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17] = !N14562;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0] = (N11888 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[17]) | ((!N11888) & N11890);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38 = float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 = !((float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__34) | float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__33);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[7]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[6]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[5]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[4]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[3]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[2]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[1]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23] = (float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42 & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__22[0]) | ((!float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__42) & float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__38);
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31] = !(float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__29 | (!a_sign));
reg x_reg_L0_23__I2278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__I2278_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[23];
	end
assign N5677 = x_reg_L0_23__I2278_QOUT;
reg x_reg_L0_24__I2279_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_24__I2279_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[24];
	end
assign N5682 = x_reg_L0_24__I2279_QOUT;
reg x_reg_L0_25__I2280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_25__I2280_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[25];
	end
assign N5687 = x_reg_L0_25__I2280_QOUT;
reg x_reg_L0_26__I2281_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_26__I2281_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[26];
	end
assign N5692 = x_reg_L0_26__I2281_QOUT;
reg x_reg_L0_27__I2282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_27__I2282_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[27];
	end
assign N5697 = x_reg_L0_27__I2282_QOUT;
reg x_reg_L0_28__I2283_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_28__I2283_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[28];
	end
assign N5702 = x_reg_L0_28__I2283_QOUT;
reg x_reg_L0_29__I2284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__I2284_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[29];
	end
assign N5707 = x_reg_L0_29__I2284_QOUT;
reg x_reg_L0_30__I2285_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_30__I2285_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[30];
	end
assign N5712 = x_reg_L0_30__I2285_QOUT;
reg x_reg_L0_31__I2286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I2286_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[31];
	end
assign N5717 = x_reg_L0_31__I2286_QOUT;
reg x_reg_L1_0__I2287_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__I2287_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[0];
	end
assign x[0] = x_reg_L1_0__I2287_QOUT;
reg x_reg_L1_1__I2288_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__I2288_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[1];
	end
assign x[1] = x_reg_L1_1__I2288_QOUT;
reg x_reg_L1_2__I2289_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__I2289_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[2];
	end
assign x[2] = x_reg_L1_2__I2289_QOUT;
reg x_reg_L1_3__I2290_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__I2290_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[3];
	end
assign x[3] = x_reg_L1_3__I2290_QOUT;
reg x_reg_L1_4__I2291_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__I2291_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[4];
	end
assign x[4] = x_reg_L1_4__I2291_QOUT;
reg x_reg_L1_5__I2292_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__I2292_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[5];
	end
assign x[5] = x_reg_L1_5__I2292_QOUT;
reg x_reg_L1_6__I2293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__I2293_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[6];
	end
assign x[6] = x_reg_L1_6__I2293_QOUT;
reg x_reg_L1_7__I2294_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__I2294_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[7];
	end
assign x[7] = x_reg_L1_7__I2294_QOUT;
reg x_reg_L1_8__I2295_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__I2295_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[8];
	end
assign x[8] = x_reg_L1_8__I2295_QOUT;
reg x_reg_L1_9__I2296_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__I2296_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[9];
	end
assign x[9] = x_reg_L1_9__I2296_QOUT;
reg x_reg_L1_10__I2297_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__I2297_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[10];
	end
assign x[10] = x_reg_L1_10__I2297_QOUT;
reg x_reg_L1_11__I2298_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__I2298_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[11];
	end
assign x[11] = x_reg_L1_11__I2298_QOUT;
reg x_reg_L1_12__I2299_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__I2299_QOUT <= float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[12];
	end
assign x[12] = x_reg_L1_12__I2299_QOUT;
reg x_reg_L1_23__I2310_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__I2310_QOUT <= N5677;
	end
assign x[23] = x_reg_L1_23__I2310_QOUT;
reg x_reg_L1_24__I2311_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_24__I2311_QOUT <= N5682;
	end
assign x[24] = x_reg_L1_24__I2311_QOUT;
reg x_reg_L1_25__I2312_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_25__I2312_QOUT <= N5687;
	end
assign x[25] = x_reg_L1_25__I2312_QOUT;
reg x_reg_L1_26__I2313_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_26__I2313_QOUT <= N5692;
	end
assign x[26] = x_reg_L1_26__I2313_QOUT;
reg x_reg_L1_27__I2314_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_27__I2314_QOUT <= N5697;
	end
assign x[27] = x_reg_L1_27__I2314_QOUT;
reg x_reg_L1_28__I2315_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_28__I2315_QOUT <= N5702;
	end
assign x[28] = x_reg_L1_28__I2315_QOUT;
reg x_reg_L1_29__I2316_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__I2316_QOUT <= N5707;
	end
assign x[29] = x_reg_L1_29__I2316_QOUT;
reg x_reg_L1_30__I2317_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_30__I2317_QOUT <= N5712;
	end
assign x[30] = x_reg_L1_30__I2317_QOUT;
reg x_reg_L1_31__I2318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I2318_QOUT <= N5717;
	end
assign x[31] = x_reg_L1_31__I2318_QOUT;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[14] = x[14];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[15] = x[15];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[16] = x[16];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[17] = x[17];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[18] = x[18];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[19] = x[19];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[20] = x[20];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[21] = x[21];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[22] = x[22];
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_x[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__19[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__20[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__51[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[16] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[17] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[18] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[19] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__60[20] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[25] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[26] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[27] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[28] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[29] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[30] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[31] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[32] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[33] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__62__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W0[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[34] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[35] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[36] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[37] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[38] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__63__W1[39] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[0] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[1] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[2] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[3] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[4] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[5] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[6] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[7] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[8] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[9] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[10] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[11] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[12] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[13] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[14] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[15] = 1'B0;
assign float_div_cynw_cm_float_rcp_E8_M23_3_inst_inst_cellmath__64[16] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  vLf3SQnarR8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



