/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:20 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_2_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__4,
	inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49,
	inst_cellmath__51;
wire N440,N441,N442,N444,N445,N446,N447 
	,N450,N461,N469,N470,N1900,N1902,N1923,N1931 
	,N1934,N1936,N1940,N1942,N1945,N1951,N1955,N1980 
	,N1985,N1989,N1992,N2011,N2013,N2034,N2042,N2045 
	,N2047,N2051,N2053,N2056,N2062,N2066,N2091,N2096 
	,N2100,N2103,N2135,N2140,N2147,N2148,N2149,N2150 
	,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158 
	,N2159,N2160,N2161,N2162,N2163,N2164,N2166,N2167 
	,N2168,N2169,N2170,N2171,N2172,N2173,N2174,N2175 
	,N2177,N2178,N2179,N2180,N2181,N2183,N2184,N2185 
	,N2186,N2187,N2188,N2189,N2190,N2191,N2192,N2193 
	,N2194,N2195,N2196,N2197,N2198,N2199,N2200,N2201 
	,N2202,N2203,N2204,N2205,N2206,N2207,N2208,N2209 
	,N2210,N2211,N2212,N2213,N2214,N2215,N2216,N2217 
	,N2218,N2219,N2220,N2221,N2222,N2224,N2225,N2227 
	,N2228,N2229,N2230,N2231,N2232,N2233,N2234,N2235 
	,N2236,N2237,N2238,N2241,N2242,N2243,N2244,N2245 
	,N2247,N2248,N2249,N2250,N2251,N2252,N2253,N2254 
	,N2255,N2256,N2257,N2258,N2259,N2260,N2261,N2262 
	,N2263,N2264,N2265,N2266,N2267,N2268,N2269,N2270 
	,N2271,N2272,N2273,N2274,N2275,N2276,N2277,N2278 
	,N2279,N2281,N2282,N2283,N2284,N2285,N2286,N2287 
	,N2288,N2289,N2290,N2291,N2292,N2293,N2294,N2295 
	,N2296,N2297,N2298,N2299,N2300,N2302,N2303,N2305 
	,N2306,N2307,N2308,N2309,N2310,N2311,N2312,N2313 
	,N2314,N2315,N2316,N2317,N2318,N2319,N2320,N2321 
	,N2322,N2323,N2325,N2326,N2327,N2328,N2329,N2330 
	,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338 
	,N2339,N2340,N2341,N2343,N2344,N2345,N2346,N2347 
	,N2348,N2349,N2350,N2351,N2352,N2353,N2354,N2355 
	,N2356,N2357,N2358,N2359,N2360,N2361,N2362,N2363 
	,N2364,N2366,N2367,N2368,N2370,N2371,N2372,N2373 
	,N2374,N2375,N2376,N2377,N2378,N2379,N2381,N2382 
	,N2383,N2384,N2385,N2386,N2387,N2389,N2390,N2391 
	,N2392,N2393,N2394,N2395,N2396,N2397,N2398,N2399 
	,N2400,N2401,N2402,N2403,N2404,N2405,N2406,N2407 
	,N2408,N2409,N2410,N2411,N2412,N2413,N2414,N2415 
	,N2416,N2417,N2418,N2420,N2421,N2423,N2424,N2425 
	,N2426,N2427,N2428,N2429,N2430,N2431,N2432,N2433 
	,N2435,N2436,N2437,N2438,N2439,N2440,N2441,N2442 
	,N2443,N2445,N2446,N2447,N2448,N2449,N2450,N2451 
	,N2452,N2453,N2454,N2455,N2456,N2457,N2458,N2459 
	,N2460,N2461,N2462,N2463,N2465,N2466,N2467,N2468 
	,N2469,N2470,N2471,N2472,N2473,N2474,N2475,N2476 
	,N2478,N2479,N2480,N2481,N2482,N2483,N2484,N2485 
	,N2486,N2487,N2488,N2489,N2490,N2491,N2492,N2493 
	,N2494,N2495,N2496,N2497,N2498,N2499,N2501,N2502 
	,N2503,N2504,N2506,N2507,N2508,N2509,N2511,N2512 
	,N2513,N2514,N2515,N2516,N2517,N2518,N2519,N2520 
	,N2521,N2522,N2523,N2525,N2526,N2527,N2528,N2529 
	,N2530,N2531,N2532,N2533,N2534,N2535,N2536,N2537 
	,N2538,N2539,N2540,N2541,N2542,N2543,N2544,N2545 
	,N2546,N2547,N2548,N2549,N2550,N2551,N2552,N2553 
	,N2554,N2555,N2556,N2557,N2558,N2559,N2560,N2561 
	,N2562,N2563,N2564,N2566,N2567,N2568,N2570,N2571 
	,N2572,N2573,N2574,N2575,N2576,N2577,N2578,N2579 
	,N2580,N2581,N2582,N2583,N2584,N2585,N2586,N2588 
	,N2589,N2590,N2591,N2592,N2594,N2595,N2596,N2597 
	,N2598,N2599,N2600,N2601,N2602,N2603,N2604,N2605 
	,N2606,N2607,N2608,N2609,N2610,N2611,N2612,N2613 
	,N2614,N2615,N2616,N2617,N2618,N2620,N2621,N2622 
	,N2623,N2624,N2625,N2626,N2628,N2629,N2630,N2631 
	,N2633,N2634,N2635,N2636,N2637,N2638,N2639,N2640 
	,N2641,N2642,N2643,N2644,N2645,N2646,N2648,N2649 
	,N2650,N2651,N2652,N2653,N2654,N2655,N2656,N2657 
	,N2658,N2659,N2660,N2661,N2662,N2663,N2664,N2666 
	,N2667,N2668,N2669,N2670,N2671,N2672,N2673,N2674 
	,N2675,N2676,N2677,N2678,N2679,N2680,N2682,N2683 
	,N2684,N2685,N2686,N2687,N2688,N2689,N2690,N2691 
	,N2692,N2693,N2694,N2695,N2696,N2697,N2698,N2699 
	,N2700,N2701,N2702,N2703,N2704,N2705,N2706,N2708 
	,N2709,N2710,N2712,N2713,N2714,N2715,N2716,N2717 
	,N2718,N2719,N2720,N2721,N2723,N2724,N2725,N2726 
	,N2727,N2728,N2729,N2730,N2731,N2732,N2733,N2734 
	,N2735,N2736,N2737,N2738,N2739,N2740,N2741,N2742 
	,N2743,N2744,N2745,N2746,N2747,N2748,N2749,N2750 
	,N2751,N2752,N2753,N2754,N2755,N2756,N2757,N2758 
	,N2759,N2760,N2761,N2762,N2763,N2764,N2765,N2767 
	,N2768,N2769,N2770,N2771,N2772,N2773,N2774,N2775 
	,N2776,N2777,N2778,N2779,N2780,N2781,N2782,N2783 
	,N2785,N2786,N2787,N2788,N2789,N2790,N2791,N2793 
	,N2794,N2795,N2796,N2797,N2798,N2799,N2800,N2801 
	,N2802,N2803,N2804,N2805,N2806,N2807,N2808,N2809 
	,N2810,N2811,N2812,N2813,N2814,N2815,N2816,N2817 
	,N2818,N2819,N2820,N2821,N2822,N2824,N2825,N2826 
	,N2827,N2828,N2829,N2831,N2832,N2833,N2834,N2835 
	,N2836,N2837,N2838,N2839,N2840,N2841,N2842,N2843 
	,N2844,N2845,N2846,N2847,N2849,N2850,N2851,N2852 
	,N2853,N2854,N2855,N2856,N2857,N2858,N2859,N2860 
	,N2861,N2862,N2863,N2864,N2865,N2867,N2868,N2869 
	,N2870,N2871,N2872,N2873,N2874,N2875,N2876,N2877 
	,N2878,N2879,N2880,N2881,N2882,N2883,N2884,N2885 
	,N2886,N2887,N2888,N2889,N2890,N2891,N2892,N2893 
	,N2894,N2895,N2896,N2897,N2898,N2899,N2900,N2901 
	,N2902,N2903,N2905,N2906,N2908,N2909,N2910,N2911 
	,N2912,N2913,N2914,N2915,N2916,N2917,N2918,N2919 
	,N2920,N2922,N2923,N2924,N2925,N2926,N2927,N2928 
	,N2929,N2931,N2932,N2933,N2934,N2935,N2936,N2937 
	,N2938,N2939,N2940,N2941,N2942,N2943,N2944,N2945 
	,N2946,N2947,N2948,N2949,N2950,N2951,N2952,N2953 
	,N2954,N2955,N2956,N2957,N2959,N2960,N2961,N2962 
	,N2963,N2964,N2965,N2966,N2967,N2968,N2969,N2970 
	,N2971,N2972,N2973,N2974,N2975,N2976,N2977,N2978 
	,N2979,N2980,N2981,N2983,N2984,N2985,N2986,N2987 
	,N2988,N2989,N2990,N2991,N2992,N2993,N2994,N2995 
	,N2996,N2997,N2998,N2999,N3001,N3002,N3003,N3004 
	,N3005,N3006,N3007,N3008,N3009,N3010,N3011,N3012 
	,N3013,N3014,N3015,N3016,N3018,N3019,N3020,N3021 
	,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029 
	,N3030,N3031,N3032,N3033,N3034,N3035,N3036,N3037 
	,N3038,N3039,N3040,N3041,N3042,N3044,N3045,N3046 
	,N3047,N3048,N3049,N3050,N3051,N3052,N3053,N3054 
	,N3055,N3056,N3057,N3058,N3060,N3061,N3062,N3063 
	,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071 
	,N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079 
	,N3080,N3081,N3082,N3083,N3084,N3085,N3086,N3087 
	,N3088,N3089,N3090,N3091,N3092,N3093,N3094,N3095 
	,N3096,N3097,N3098,N3099,N3100,N3102,N3103,N3104 
	,N3105,N3106,N3107,N3109,N3110,N3111,N3112,N3113 
	,N3114,N3115,N3116,N3117,N3118,N3119,N3121,N3122 
	,N3123,N3124,N3125,N3126,N3128,N3129,N3130,N3131 
	,N3132,N3133,N3134,N3135,N3136,N3137,N3138,N3139 
	,N3140,N3141,N3142,N3143,N3144,N3145,N3146,N3147 
	,N3148,N3149,N3150,N3151,N3152,N3153,N3154,N3155 
	,N3156,N3158,N3159,N3160,N3161,N3162,N3163,N3164 
	,N3165,N3166,N3167,N3168,N3169,N3170,N3171,N3172 
	,N3173,N3174,N3175,N3176,N3177,N3178,N3179,N3182 
	,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190 
	,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3199 
	,N3200,N3201,N3202,N3203,N3204,N3205,N3206,N3207 
	,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215 
	,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223 
	,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231 
	,N3232,N3233,N3234,N3235,N3236,N3237,N3239,N3240 
	,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248 
	,N3249,N3250,N3251,N3252,N3253,N3254,N3255,N3256 
	,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265 
	,N3267,N3268,N3269,N3270,N3271,N3272,N3273,N3274 
	,N3275,N3276,N3277,N3278,N3279,N3280,N3281,N3282 
	,N3283,N3284,N3285,N3286,N3287,N3288,N3289,N3290 
	,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3299 
	,N3300,N3302,N3303,N3304,N3305,N3306,N3307,N3308 
	,N3309,N3310,N3311,N3312,N3313,N3314,N3315,N3316 
	,N3317,N3318,N3319,N3320,N3321,N3323,N3324,N3325 
	,N3326,N3327,N3328,N3329,N3330,N3331,N3332,N3333 
	,N3334,N3335,N3336,N3337,N3338,N3339,N3340,N3341 
	,N3342,N3344,N3345,N3346,N3347,N3348,N3349,N3350 
	,N3351,N3352,N3353,N3354,N3355,N3356,N3357,N3358 
	,N3360,N3361,N3362,N3363,N3364,N3365,N3366,N3367 
	,N3368,N3369,N3370,N3371,N3372,N3373,N3374,N3375 
	,N3376,N3377,N3379,N3380,N3381,N3384,N3385,N3386 
	,N3388,N3389,N3390,N3391,N3392,N3393,N3394,N3395 
	,N3396,N3397,N3398,N3399,N3400,N3401,N3402,N3403 
	,N3405,N3406,N3407,N3408,N3409,N3410,N3411,N3412 
	,N3413,N3414,N3415,N3416,N3417,N3418,N3419,N3420 
	,N3421,N3422,N3423,N3424,N3425,N3426,N3427,N3428 
	,N3429,N3430,N3431,N3432,N3433,N3434,N3435,N3436 
	,N3437,N3438,N3439,N3441,N3442,N3443,N3444,N3445 
	,N3446,N3447,N3448,N3449,N3450,N3451,N3452,N3454 
	,N3455,N3456,N3457,N3458,N3459,N3460,N3462,N3463 
	,N3464,N3465,N3466,N3467,N3468,N3469,N3470,N3471 
	,N3472,N3473,N3474,N3475,N3476,N3477,N3478,N3479 
	,N3480,N3481,N3482,N3483,N3484,N3485,N3487,N3488 
	,N3489,N3491,N3492,N3493,N3494,N3495,N3496,N3497 
	,N3498,N3499,N3500,N3501,N3502,N3503,N3504,N3505 
	,N3506,N3507,N3508,N3510,N3511,N3512,N3513,N3514 
	,N3515,N3516,N3517,N3518,N3519,N3520,N3521,N3522 
	,N3523,N3524,N3525,N3526,N3527,N3528,N3530,N3531 
	,N3532,N3533,N3534,N3535,N3536,N3537,N3538,N3539 
	,N3540,N3541,N3542,N3544,N3545,N3546,N3547,N3548 
	,N3549,N3550,N3551,N3552,N3553,N3554,N3555,N3556 
	,N3557,N3558,N3560,N3561,N3562,N3563,N3564,N3565 
	,N3566,N3567,N3568,N3569,N3570,N3571,N3573,N3574 
	,N3575,N3576,N3578,N3579,N3580,N3581,N3582,N3583 
	,N3584,N3585,N3586,N3587,N3588,N3589,N3590,N3592 
	,N3593,N3594,N3596,N3597,N3599,N3600,N3601,N3602 
	,N3603,N3604,N3605,N3606,N3607,N3608,N3609,N3610 
	,N3611,N3612,N3613,N3614,N3615,N3616,N3617,N3618 
	,N3619,N3620,N3621,N3622,N3623,N3624,N3625,N3626 
	,N3627,N3628,N3629,N3630,N3632,N3633,N3634,N3635 
	,N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643 
	,N3644,N3645,N3646,N3647,N3648,N3649,N3650,N3651 
	,N3652,N3654,N3655,N3656,N3658,N3659,N3660,N3661 
	,N3662,N3663,N3664,N3665,N3666,N3667,N3668,N3669 
	,N3670,N3672,N3673,N3674,N3675,N3676,N3677,N3678 
	,N3679,N3680,N3681,N3682,N3683,N3684,N3686,N3687 
	,N3688,N3689,N5224,N5333,N5336,N5337,N5338,N5341 
	,N5344,N5345,N5346,N5351,N5353,N5359,N5361,N5363 
	,N5365,N5366,N5369,N5370,N5371,N5373,N5375,N5378 
	,N5384,N5385,N5387,N5390,N5392,N5394,N5400,N5403 
	,N5404,N5405,N5406,N5408,N5411,N5412,N5416,N5419 
	,N5422,N5500,N5528,N5530,N5532,N5536,N5538,N5540 
	,N5543,N5545,N5547,N5552,N5554,N5558,N5624,N5627 
	,N5631,N5632,N5637,N5643,N5647,N5652,N5655,N5681 
	,N5682,N5690,N5691,N5697,N5699,N5700,N5701,N5763 
	,N5768,N5772,N5775,N5801,N5808,N5812,N5813,N5815 
	,N5823,N5830,N5852,N5860,N5870,N5874,N5884,N5887 
	,N5893,N5914,N5923,N5925,N5930,N5931,N5933,N5934 
	,N5941,N5943,N5948,N5951,N5953,N5955,N5957,N5959 
	,N5965,N5967,N5970,N5973,N5977,N5978,N5980,N5982 
	,N5984,N5987,N5990,N5992,N5996,N5999,N6002,N6004 
	,N6005,N6008,N6014,N6016,N6018,N6020,N6024,N6027 
	,N6028,N6030,N6032,N6038,N6040,N6043,N6047,N6048 
	,N6051,N6053,N6055,N6061,N6063,N6066,N6069,N6073 
	,N6075,N6077,N6079,N6080,N6084,N6086,N6088,N6091 
	,N6095,N6096,N6098,N6100,N6102,N6104,N6109,N6112 
	,N6114,N6117,N8295,N8298,N8302,N8310,N8320,N8325 
	,N8327,N8328,N8334,N8335,N8336,N8342,N8343,N8352 
	,N8358,N8359,N8368,N8373,N8376,N8378,N8380,N8382 
	,N8388,N8396,N8402,N8411,N8417;
NAND2XL inst_cellmath__17_0_I272 (.Y(N1900), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__17_0_I10192 (.Y(N1902), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3706 (.Y(N8388), .A(b_exp[7]), .B(b_exp[6]), .C(N1902));
NOR2XL hyperpropagate_4_1_A_I3707 (.Y(inst_cellmath__17), .A(N1900), .B(N8388));
NOR2XL inst_cellmath__19__2__I285 (.Y(N1923), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__19__2__I286 (.Y(N1931), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__19__2__I287 (.Y(N1942), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__19__2__I288 (.Y(N1951), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__19__2__I10193 (.Y(N1936), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__19__2__I10194 (.Y(N1945), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__19__2__I10195 (.Y(N1955), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__19__2__I292 (.Y(N1940), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N1936));
NAND4XL inst_cellmath__19__2__I294 (.Y(N1934), .A(N1923), .B(N1942), .C(N1931), .D(N1951));
NOR4BX1 inst_cellmath__19__2__I10196 (.Y(inst_cellmath__19), .AN(N1940), .B(N1934), .C(N1945), .D(N1955));
NAND2XL cynw_cm_float_mul_ieee_I297 (.Y(inst_cellmath__21), .A(inst_cellmath__17), .B(inst_cellmath__19));
NOR2XL inst_cellmath__13__1__I298 (.Y(N1985), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL inst_cellmath__13__1__I299 (.Y(N1989), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__13__1__I300 (.Y(N1992), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__13__1__I301 (.Y(N1980), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__13__1__I3679 (.Y(inst_cellmath__13), .A(N1985), .B(N1992), .C(N1989), .D(N1980));
NOR2XL cynw_cm_float_mul_ieee_I305 (.Y(N441), .A(inst_cellmath__13), .B(inst_cellmath__21));
NAND2XL inst_cellmath__10_0_I306 (.Y(N2011), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__10_0_I10197 (.Y(N2013), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3708 (.Y(N8396), .A(a_exp[7]), .B(a_exp[6]), .C(N2013));
NOR2XL hyperpropagate_4_1_A_I3709 (.Y(inst_cellmath__10), .A(N2011), .B(N8396));
NOR2XL inst_cellmath__12__0__I319 (.Y(N2034), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__12__0__I320 (.Y(N2042), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__12__0__I321 (.Y(N2053), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__12__0__I322 (.Y(N2062), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__12__0__I10198 (.Y(N2047), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__12__0__I10199 (.Y(N2056), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__12__0__I10200 (.Y(N2066), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__12__0__I326 (.Y(N2051), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N2047));
NAND4XL inst_cellmath__12__0__I328 (.Y(N2045), .A(N2034), .B(N2053), .C(N2042), .D(N2062));
NOR4BX1 inst_cellmath__12__0__I10201 (.Y(inst_cellmath__12), .AN(N2051), .B(N2045), .C(N2056), .D(N2066));
NAND2XL cynw_cm_float_mul_ieee_I331 (.Y(inst_cellmath__14), .A(inst_cellmath__10), .B(inst_cellmath__12));
NOR2XL inst_cellmath__20__3__I332 (.Y(N2096), .A(b_exp[0]), .B(b_exp[1]));
NOR2XL inst_cellmath__20__3__I333 (.Y(N2100), .A(b_exp[7]), .B(b_exp[6]));
NOR2XL inst_cellmath__20__3__I334 (.Y(N2103), .A(b_exp[5]), .B(b_exp[4]));
NOR2XL inst_cellmath__20__3__I335 (.Y(N2091), .A(b_exp[3]), .B(b_exp[2]));
NAND4XL inst_cellmath__20__3__I3681 (.Y(inst_cellmath__20), .A(N2096), .B(N2103), .C(N2100), .D(N2091));
NOR2XL cynw_cm_float_mul_ieee_I339 (.Y(N440), .A(inst_cellmath__20), .B(inst_cellmath__14));
NOR2BX1 cynw_cm_float_mul_ieee_I340 (.Y(inst_cellmath__15), .AN(inst_cellmath__10), .B(inst_cellmath__12));
NOR2BX1 cynw_cm_float_mul_ieee_I341 (.Y(inst_cellmath__22), .AN(inst_cellmath__17), .B(inst_cellmath__19));
OR4X1 cynw_cm_float_mul_ieee_I342 (.Y(inst_cellmath__26), .A(inst_cellmath__22), .B(inst_cellmath__15), .C(N441), .D(N440));
XOR2XL cynw_cm_float_mul_ieee_I343 (.Y(inst_cellmath__23), .A(a_sign), .B(b_sign));
NAND2BXL inst_cellmath__41_0_I344 (.Y(N2135), .AN(b_sign), .B(inst_cellmath__22));
MX2XL inst_cellmath__41_0_I345 (.Y(N2140), .A(N2135), .B(a_sign), .S0(inst_cellmath__15));
MX2XL inst_cellmath__41_0_I346 (.Y(x[31]), .A(inst_cellmath__23), .B(N2140), .S0(inst_cellmath__26));
INVXL inst_cellmath__24_0_I347 (.Y(N3445), .A(a_man[0]));
INVXL inst_cellmath__24_0_I348 (.Y(N2228), .A(a_man[1]));
INVXL inst_cellmath__24_0_I349 (.Y(N2573), .A(a_man[2]));
INVXL inst_cellmath__24_0_I350 (.Y(N2911), .A(a_man[3]));
INVXL inst_cellmath__24_0_I351 (.Y(N3243), .A(a_man[4]));
INVXL inst_cellmath__24_0_I352 (.Y(N3578), .A(a_man[5]));
INVXL inst_cellmath__24_0_I353 (.Y(N2368), .A(a_man[6]));
INVXL inst_cellmath__24_0_I354 (.Y(N2713), .A(a_man[7]));
INVXL inst_cellmath__24_0_I355 (.Y(N3047), .A(a_man[8]));
INVXL inst_cellmath__24_0_I356 (.Y(N3391), .A(a_man[9]));
INVXL inst_cellmath__24_0_I357 (.Y(N2171), .A(a_man[10]));
INVXL inst_cellmath__24_0_I358 (.Y(N2511), .A(a_man[11]));
INVXL inst_cellmath__24_0_I359 (.Y(N2853), .A(a_man[12]));
INVXL inst_cellmath__24_0_I360 (.Y(N3186), .A(a_man[13]));
INVXL inst_cellmath__24_0_I361 (.Y(N3513), .A(a_man[14]));
INVXL inst_cellmath__24_0_I362 (.Y(N2308), .A(a_man[15]));
INVXL inst_cellmath__24_0_I363 (.Y(N2653), .A(a_man[16]));
INVXL inst_cellmath__24_0_I364 (.Y(N2987), .A(a_man[17]));
INVXL inst_cellmath__24_0_I365 (.Y(N3329), .A(a_man[18]));
INVXL inst_cellmath__24_0_I366 (.Y(N3660), .A(a_man[19]));
INVXL inst_cellmath__24_0_I367 (.Y(N2452), .A(a_man[20]));
INVXL inst_cellmath__24_0_I368 (.Y(N2799), .A(a_man[21]));
INVXL inst_cellmath__24_0_I369 (.Y(N3134), .A(a_man[22]));
INVXL inst_cellmath__24_0_I370 (.Y(N2357), .A(b_man[0]));
NAND2X2 inst_cellmath__24_0_I371 (.Y(N2935), .A(b_man[1]), .B(N2357));
INVX1 inst_cellmath__24_0_I372 (.Y(N3272), .A(b_man[1]));
XNOR2X1 inst_cellmath__24_0_I373 (.Y(N2636), .A(N3445), .B(N3272));
OAI22XL inst_cellmath__24_0_I374 (.Y(N2292), .A0(N2636), .A1(N2357), .B0(N3272), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I375 (.Y(N3312), .A(N2228), .B(N3272));
OAI22XL inst_cellmath__24_0_I376 (.Y(N2217), .A0(N3312), .A1(N2357), .B0(N2636), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I377 (.Y(N2437), .A(N2573), .B(N3272));
OAI22XL inst_cellmath__24_0_I378 (.Y(N3647), .A0(N2437), .A1(N2357), .B0(N3312), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I379 (.Y(N3116), .A(N2911), .B(N3272));
OAI22XL inst_cellmath__24_0_I380 (.Y(N2781), .A0(N3116), .A1(N2357), .B0(N2437), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I381 (.Y(N2237), .A(N3243), .B(N3272));
OAI22XL inst_cellmath__24_0_I382 (.Y(N3452), .A0(N2237), .A1(N2357), .B0(N3116), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I383 (.Y(N2920), .A(N3578), .B(N3272));
OAI22XL inst_cellmath__24_0_I384 (.Y(N2584), .A0(N2920), .A1(N2357), .B0(N2237), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I385 (.Y(N3588), .A(N2368), .B(N3272));
OAI22XL inst_cellmath__24_0_I386 (.Y(N3253), .A0(N3588), .A1(N2357), .B0(N2920), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I387 (.Y(N2720), .A(N2713), .B(N3272));
OAI22XL inst_cellmath__24_0_I388 (.Y(N2378), .A0(N2720), .A1(N2357), .B0(N3588), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I389 (.Y(N3401), .A(N3047), .B(N3272));
OAI22XL inst_cellmath__24_0_I390 (.Y(N3054), .A0(N3401), .A1(N2357), .B0(N2720), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I391 (.Y(N2521), .A(N3391), .B(N3272));
OAI22XL inst_cellmath__24_0_I392 (.Y(N2180), .A0(N2521), .A1(N2357), .B0(N3401), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I393 (.Y(N3195), .A(N2171), .B(N3272));
OAI22XL inst_cellmath__24_0_I394 (.Y(N2863), .A0(N3195), .A1(N2357), .B0(N2521), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I395 (.Y(N2321), .A(N2511), .B(N3272));
OAI22XL inst_cellmath__24_0_I396 (.Y(N3525), .A0(N2321), .A1(N2357), .B0(N3195), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I397 (.Y(N2998), .A(N2853), .B(N3272));
OAI22XL inst_cellmath__24_0_I398 (.Y(N2664), .A0(N2998), .A1(N2357), .B0(N2321), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I399 (.Y(N3669), .A(N3186), .B(N3272));
OAI22XL inst_cellmath__24_0_I400 (.Y(N3341), .A0(N3669), .A1(N2357), .B0(N2998), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I401 (.Y(N2808), .A(N3513), .B(N3272));
OAI22XL inst_cellmath__24_0_I402 (.Y(N2461), .A0(N2808), .A1(N2357), .B0(N3669), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I403 (.Y(N3471), .A(N2308), .B(N3272));
OAI22XL inst_cellmath__24_0_I404 (.Y(N3143), .A0(N3471), .A1(N2357), .B0(N2808), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I405 (.Y(N2604), .A(N2653), .B(N3272));
OAI22XL inst_cellmath__24_0_I406 (.Y(N2263), .A0(N2604), .A1(N2357), .B0(N3471), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I407 (.Y(N3280), .A(N2987), .B(N3272));
OAI22XL inst_cellmath__24_0_I408 (.Y(N2943), .A0(N3280), .A1(N2357), .B0(N2604), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I409 (.Y(N2401), .A(N3329), .B(N3272));
OAI22XL inst_cellmath__24_0_I410 (.Y(N3615), .A0(N2401), .A1(N2357), .B0(N3280), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I411 (.Y(N3083), .A(N3660), .B(N3272));
OAI22XL inst_cellmath__24_0_I412 (.Y(N2749), .A0(N3083), .A1(N2357), .B0(N2401), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I413 (.Y(N2204), .A(N2452), .B(N3272));
OAI22XL inst_cellmath__24_0_I414 (.Y(N3424), .A0(N2204), .A1(N2357), .B0(N3083), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I415 (.Y(N2888), .A(N2799), .B(N3272));
OAI22XL inst_cellmath__24_0_I416 (.Y(N2548), .A0(N2888), .A1(N2357), .B0(N2204), .B1(N2935));
XNOR2X1 inst_cellmath__24_0_I417 (.Y(N3553), .A(N3134), .B(N3272));
OAI22XL inst_cellmath__24_0_I418 (.Y(N3221), .A0(N3553), .A1(N2357), .B0(N2888), .B1(N2935));
INVXL inst_cellmath__24_0_I419 (.Y(N2691), .A(N3272));
OAI22XL inst_cellmath__24_0_I420 (.Y(N2350), .A0(N2691), .A1(N2357), .B0(N3553), .B1(N2935));
MXI2XL inst_cellmath__24_0_I421 (.Y(N3024), .A(N2935), .B(N2357), .S0(N2691));
XNOR2X1 inst_cellmath__24_0_I422 (.Y(N2968), .A(b_man[2]), .B(b_man[1]));
INVXL inst_cellmath__24_0_I3558 (.Y(N8295), .A(N2968));
INVXL inst_cellmath__24_0_I3565 (.Y(N8302), .A(N8295));
INVXL inst_cellmath__24_0_I3561 (.Y(N8298), .A(N8295));
XOR2XL inst_cellmath__24_0_I423 (.Y(N2211), .A(b_man[3]), .B(b_man[1]));
NAND2X2 inst_cellmath__24_0_I424 (.Y(N2620), .A(N2211), .B(N2968));
INVX1 inst_cellmath__24_0_I425 (.Y(N2959), .A(b_man[3]));
NAND2XL inst_cellmath__24_0_I426 (.Y(N3111), .A(b_man[1]), .B(b_man[2]));
AND2XL inst_cellmath__24_0_I427 (.Y(N3446), .A(b_man[3]), .B(N3111));
XNOR2X1 inst_cellmath__24_0_I428 (.Y(N2577), .A(N3445), .B(N2959));
OAI22XL inst_cellmath__24_0_I429 (.Y(N2231), .A0(N2577), .A1(N8302), .B0(N2959), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I430 (.Y(N3246), .A(N2228), .B(N2959));
OAI22XL inst_cellmath__24_0_I431 (.Y(N2913), .A0(N3246), .A1(N8302), .B0(N2577), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I432 (.Y(N2370), .A(N2573), .B(N2959));
OAI22XL inst_cellmath__24_0_I433 (.Y(N3582), .A0(N2370), .A1(N8302), .B0(N3246), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I434 (.Y(N3051), .A(N2911), .B(N2959));
OAI22XL inst_cellmath__24_0_I435 (.Y(N2715), .A0(N3051), .A1(N8302), .B0(N2370), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I436 (.Y(N2173), .A(N3243), .B(N2959));
OAI22XL inst_cellmath__24_0_I437 (.Y(N3396), .A0(N2173), .A1(N8302), .B0(N3051), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I438 (.Y(N2858), .A(N3578), .B(N2959));
OAI22XL inst_cellmath__24_0_I439 (.Y(N2517), .A0(N2858), .A1(N8302), .B0(N2173), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I440 (.Y(N3519), .A(N2368), .B(N2959));
OAI22XL inst_cellmath__24_0_I441 (.Y(N3188), .A0(N3519), .A1(N8302), .B0(N2858), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I442 (.Y(N2655), .A(N2713), .B(N2959));
OAI22XL inst_cellmath__24_0_I443 (.Y(N2314), .A0(N2655), .A1(N8302), .B0(N3519), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I444 (.Y(N3334), .A(N3047), .B(N2959));
OAI22XL inst_cellmath__24_0_I445 (.Y(N2991), .A0(N3334), .A1(N8302), .B0(N2655), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I446 (.Y(N2455), .A(N3391), .B(N2959));
OAI22XL inst_cellmath__24_0_I447 (.Y(N3662), .A0(N2455), .A1(N8302), .B0(N3334), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I448 (.Y(N3135), .A(N2171), .B(N2959));
OAI22XL inst_cellmath__24_0_I449 (.Y(N2802), .A0(N3135), .A1(N8302), .B0(N2455), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I450 (.Y(N2257), .A(N2511), .B(N2959));
OAI22XL inst_cellmath__24_0_I451 (.Y(N3466), .A0(N2257), .A1(N8302), .B0(N3135), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I452 (.Y(N2939), .A(N2853), .B(N2959));
OAI22XL inst_cellmath__24_0_I453 (.Y(N2598), .A0(N2939), .A1(N8302), .B0(N2257), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I454 (.Y(N3608), .A(N3186), .B(N2959));
OAI22XL inst_cellmath__24_0_I455 (.Y(N3275), .A0(N3608), .A1(N8302), .B0(N2939), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I456 (.Y(N2740), .A(N3513), .B(N2959));
OAI22XL inst_cellmath__24_0_I457 (.Y(N2394), .A0(N2740), .A1(N8298), .B0(N3608), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I458 (.Y(N3417), .A(N2308), .B(N2959));
OAI22XL inst_cellmath__24_0_I459 (.Y(N3074), .A0(N3417), .A1(N8298), .B0(N2740), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I460 (.Y(N2541), .A(N2653), .B(N2959));
OAI22XL inst_cellmath__24_0_I461 (.Y(N2196), .A0(N2541), .A1(N8298), .B0(N3417), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I462 (.Y(N3215), .A(N2987), .B(N2959));
OAI22XL inst_cellmath__24_0_I463 (.Y(N2880), .A0(N3215), .A1(N8298), .B0(N2541), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I464 (.Y(N2343), .A(N3329), .B(N2959));
OAI22XL inst_cellmath__24_0_I465 (.Y(N3545), .A0(N2343), .A1(N8298), .B0(N3215), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I466 (.Y(N3019), .A(N3660), .B(N2959));
OAI22XL inst_cellmath__24_0_I467 (.Y(N2684), .A0(N3019), .A1(N8298), .B0(N2343), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I468 (.Y(N3688), .A(N2452), .B(N2959));
OAI22XL inst_cellmath__24_0_I469 (.Y(N3361), .A0(N3688), .A1(N8298), .B0(N3019), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I470 (.Y(N2825), .A(N2799), .B(N2959));
OAI22XL inst_cellmath__24_0_I471 (.Y(N2479), .A0(N2825), .A1(N8298), .B0(N3688), .B1(N2620));
XNOR2X1 inst_cellmath__24_0_I472 (.Y(N3488), .A(N3134), .B(N2959));
OAI22XL inst_cellmath__24_0_I473 (.Y(N3162), .A0(N3488), .A1(N8302), .B0(N2825), .B1(N2620));
INVXL inst_cellmath__24_0_I474 (.Y(N2624), .A(N2959));
OAI22XL inst_cellmath__24_0_I475 (.Y(N2282), .A0(N2624), .A1(N8302), .B0(N3488), .B1(N2620));
MXI2XL inst_cellmath__24_0_I476 (.Y(N2962), .A(N2620), .B(N8302), .S0(N2624));
XOR2XL inst_cellmath__24_0_I477 (.Y(N2906), .A(b_man[4]), .B(b_man[3]));
INVX1 inst_cellmath__24_0_I3573 (.Y(N8310), .A(N2906));
XNOR2X1 inst_cellmath__24_0_I478 (.Y(N3004), .A(b_man[5]), .B(b_man[3]));
OR2XL inst_cellmath__24_0_I3653 (.Y(N2302), .A(N3004), .B(N2906));
INVX1 inst_cellmath__24_0_I482 (.Y(N2645), .A(b_man[5]));
NAND2XL inst_cellmath__24_0_I483 (.Y(N3045), .A(b_man[3]), .B(b_man[4]));
AND2XL inst_cellmath__24_0_I484 (.Y(N3385), .A(b_man[5]), .B(N3045));
XNOR2X1 inst_cellmath__24_0_I485 (.Y(N2507), .A(N3445), .B(N2645));
OAI22XL inst_cellmath__24_0_I486 (.Y(N2166), .A0(N2507), .A1(N8310), .B0(N2645), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I487 (.Y(N3183), .A(N2228), .B(N2645));
OAI22XL inst_cellmath__24_0_I488 (.Y(N2850), .A0(N3183), .A1(N8310), .B0(N2507), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I489 (.Y(N2305), .A(N2573), .B(N2645));
OAI22XL inst_cellmath__24_0_I490 (.Y(N3510), .A0(N2305), .A1(N8310), .B0(N3183), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I491 (.Y(N2984), .A(N2911), .B(N2645));
OAI22XL inst_cellmath__24_0_I492 (.Y(N2649), .A0(N2984), .A1(N8310), .B0(N2305), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I493 (.Y(N3655), .A(N3243), .B(N2645));
OAI22XL inst_cellmath__24_0_I494 (.Y(N3324), .A0(N3655), .A1(N8310), .B0(N2984), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I495 (.Y(N2796), .A(N3578), .B(N2645));
OAI22XL inst_cellmath__24_0_I496 (.Y(N2448), .A0(N2796), .A1(N8310), .B0(N3655), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I497 (.Y(N3462), .A(N2368), .B(N2645));
OAI22XL inst_cellmath__24_0_I498 (.Y(N3129), .A0(N3462), .A1(N8310), .B0(N2796), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I499 (.Y(N2594), .A(N2713), .B(N2645));
OAI22XL inst_cellmath__24_0_I500 (.Y(N2249), .A0(N2594), .A1(N8310), .B0(N3462), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I501 (.Y(N3268), .A(N3047), .B(N2645));
OAI22XL inst_cellmath__24_0_I502 (.Y(N2932), .A0(N3268), .A1(N8310), .B0(N2594), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I503 (.Y(N2390), .A(N3391), .B(N2645));
OAI22XL inst_cellmath__24_0_I504 (.Y(N3600), .A0(N2390), .A1(N8310), .B0(N3268), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I505 (.Y(N3067), .A(N2171), .B(N2645));
OAI22XL inst_cellmath__24_0_I506 (.Y(N2733), .A0(N3067), .A1(N8310), .B0(N2390), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I507 (.Y(N2191), .A(N2511), .B(N2645));
OAI22XL inst_cellmath__24_0_I508 (.Y(N3411), .A0(N2191), .A1(N8310), .B0(N3067), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I509 (.Y(N2874), .A(N2853), .B(N2645));
OAI22XL inst_cellmath__24_0_I510 (.Y(N2535), .A0(N2874), .A1(N8310), .B0(N2191), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I511 (.Y(N3537), .A(N3186), .B(N2645));
OAI22XL inst_cellmath__24_0_I512 (.Y(N3207), .A0(N3537), .A1(N8310), .B0(N2874), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I513 (.Y(N2678), .A(N3513), .B(N2645));
OAI22XL inst_cellmath__24_0_I514 (.Y(N2335), .A0(N2678), .A1(N8310), .B0(N3537), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I515 (.Y(N3351), .A(N2308), .B(N2645));
OAI22XL inst_cellmath__24_0_I516 (.Y(N3010), .A0(N3351), .A1(N8310), .B0(N2678), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I517 (.Y(N2472), .A(N2653), .B(N2645));
OAI22XL inst_cellmath__24_0_I518 (.Y(N3681), .A0(N2472), .A1(N8310), .B0(N3351), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I519 (.Y(N3153), .A(N2987), .B(N2645));
OAI22XL inst_cellmath__24_0_I520 (.Y(N2818), .A0(N3153), .A1(N8310), .B0(N2472), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I521 (.Y(N2274), .A(N3329), .B(N2645));
OAI22XL inst_cellmath__24_0_I522 (.Y(N3480), .A0(N2274), .A1(N8310), .B0(N3153), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I523 (.Y(N2954), .A(N3660), .B(N2645));
OAI22XL inst_cellmath__24_0_I524 (.Y(N2616), .A0(N2954), .A1(N8310), .B0(N2274), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I525 (.Y(N3627), .A(N2452), .B(N2645));
OAI22XL inst_cellmath__24_0_I526 (.Y(N3291), .A0(N3627), .A1(N8310), .B0(N2954), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I527 (.Y(N2760), .A(N2799), .B(N2645));
OAI22XL inst_cellmath__24_0_I528 (.Y(N2411), .A0(N2760), .A1(N8310), .B0(N3627), .B1(N2302));
XNOR2X1 inst_cellmath__24_0_I529 (.Y(N3434), .A(N3134), .B(N2645));
OAI22XL inst_cellmath__24_0_I530 (.Y(N3096), .A0(N3434), .A1(N8310), .B0(N2760), .B1(N2302));
INVXL inst_cellmath__24_0_I531 (.Y(N2562), .A(N2645));
OAI22XL inst_cellmath__24_0_I532 (.Y(N2216), .A0(N2562), .A1(N8310), .B0(N3434), .B1(N2302));
MXI2XL inst_cellmath__24_0_I533 (.Y(N2897), .A(N2302), .B(N8310), .S0(N2562));
XNOR2X1 inst_cellmath__24_0_I534 (.Y(N2844), .A(b_man[6]), .B(b_man[5]));
INVXL inst_cellmath__24_0_I3583 (.Y(N8320), .A(N2844));
INVXL inst_cellmath__24_0_I3590 (.Y(N8327), .A(N8320));
INVXL inst_cellmath__24_0_I3588 (.Y(N8325), .A(N8320));
XOR2XL inst_cellmath__24_0_I535 (.Y(N2242), .A(b_man[7]), .B(b_man[5]));
NAND2X2 inst_cellmath__24_0_I536 (.Y(N3175), .A(N2242), .B(N2844));
INVX1 inst_cellmath__24_0_I537 (.Y(N2332), .A(b_man[7]));
NAND2XL inst_cellmath__24_0_I538 (.Y(N2978), .A(b_man[5]), .B(b_man[6]));
AND2XL inst_cellmath__24_0_I539 (.Y(N3317), .A(b_man[7]), .B(N2978));
XNOR2X1 inst_cellmath__24_0_I540 (.Y(N2440), .A(N3445), .B(N2332));
OAI22XL inst_cellmath__24_0_I541 (.Y(N3650), .A0(N2440), .A1(N8327), .B0(N2332), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I542 (.Y(N3122), .A(N2228), .B(N2332));
OAI22XL inst_cellmath__24_0_I543 (.Y(N2786), .A0(N3122), .A1(N8327), .B0(N2440), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I544 (.Y(N2243), .A(N2573), .B(N2332));
OAI22XL inst_cellmath__24_0_I545 (.Y(N3457), .A0(N2243), .A1(N8327), .B0(N3122), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I546 (.Y(N2927), .A(N2911), .B(N2332));
OAI22XL inst_cellmath__24_0_I547 (.Y(N2589), .A0(N2927), .A1(N8327), .B0(N2243), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I548 (.Y(N3593), .A(N3243), .B(N2332));
OAI22XL inst_cellmath__24_0_I549 (.Y(N3261), .A0(N3593), .A1(N8327), .B0(N2927), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I550 (.Y(N2725), .A(N3578), .B(N2332));
OAI22XL inst_cellmath__24_0_I551 (.Y(N2383), .A0(N2725), .A1(N8327), .B0(N3593), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I552 (.Y(N3406), .A(N2368), .B(N2332));
OAI22XL inst_cellmath__24_0_I553 (.Y(N3062), .A0(N3406), .A1(N8325), .B0(N2725), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I554 (.Y(N2526), .A(N2713), .B(N2332));
OAI22XL inst_cellmath__24_0_I555 (.Y(N2185), .A0(N2526), .A1(N8325), .B0(N3406), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I556 (.Y(N3201), .A(N3047), .B(N2332));
OAI22XL inst_cellmath__24_0_I557 (.Y(N2869), .A0(N3201), .A1(N8325), .B0(N2526), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I558 (.Y(N2328), .A(N3391), .B(N2332));
OAI22XL inst_cellmath__24_0_I559 (.Y(N3532), .A0(N2328), .A1(N8325), .B0(N3201), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I560 (.Y(N3003), .A(N2171), .B(N2332));
OAI22XL inst_cellmath__24_0_I561 (.Y(N2669), .A0(N3003), .A1(N8325), .B0(N2328), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I562 (.Y(N3673), .A(N2511), .B(N2332));
OAI22XL inst_cellmath__24_0_I563 (.Y(N3345), .A0(N3673), .A1(N8325), .B0(N3003), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I564 (.Y(N2812), .A(N2853), .B(N2332));
OAI22XL inst_cellmath__24_0_I565 (.Y(N2467), .A0(N2812), .A1(N8325), .B0(N3673), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I566 (.Y(N3474), .A(N3186), .B(N2332));
OAI22XL inst_cellmath__24_0_I567 (.Y(N3147), .A0(N3474), .A1(N8325), .B0(N2812), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I568 (.Y(N2609), .A(N3513), .B(N2332));
OAI22XL inst_cellmath__24_0_I569 (.Y(N2266), .A0(N2609), .A1(N8325), .B0(N3474), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I570 (.Y(N3284), .A(N2308), .B(N2332));
OAI22XL inst_cellmath__24_0_I571 (.Y(N2949), .A0(N3284), .A1(N8325), .B0(N2609), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I572 (.Y(N2406), .A(N2653), .B(N2332));
OAI22XL inst_cellmath__24_0_I573 (.Y(N3620), .A0(N2406), .A1(N8325), .B0(N3284), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I574 (.Y(N3089), .A(N2987), .B(N2332));
OAI22XL inst_cellmath__24_0_I575 (.Y(N2754), .A0(N3089), .A1(N8325), .B0(N2406), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I576 (.Y(N2207), .A(N3329), .B(N2332));
OAI22XL inst_cellmath__24_0_I577 (.Y(N3428), .A0(N2207), .A1(N8325), .B0(N3089), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I578 (.Y(N2892), .A(N3660), .B(N2332));
OAI22XL inst_cellmath__24_0_I579 (.Y(N2555), .A0(N2892), .A1(N8325), .B0(N2207), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I580 (.Y(N3558), .A(N2452), .B(N2332));
OAI22XL inst_cellmath__24_0_I581 (.Y(N3226), .A0(N3558), .A1(N8325), .B0(N2892), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I582 (.Y(N2695), .A(N2799), .B(N2332));
OAI22XL inst_cellmath__24_0_I583 (.Y(N2354), .A0(N2695), .A1(N8325), .B0(N3558), .B1(N3175));
XNOR2X1 inst_cellmath__24_0_I584 (.Y(N3368), .A(N3134), .B(N2332));
OAI22XL inst_cellmath__24_0_I585 (.Y(N3030), .A0(N3368), .A1(N8327), .B0(N2695), .B1(N3175));
INVXL inst_cellmath__24_0_I586 (.Y(N2493), .A(N2332));
OAI22XL inst_cellmath__24_0_I587 (.Y(N2156), .A0(N2493), .A1(N8327), .B0(N3368), .B1(N3175));
MXI2XL inst_cellmath__24_0_I588 (.Y(N2838), .A(N3175), .B(N8327), .S0(N2493));
XNOR2X1 inst_cellmath__24_0_I589 (.Y(N2779), .A(b_man[8]), .B(b_man[7]));
INVXL inst_cellmath__24_0_I3591 (.Y(N8328), .A(N2779));
INVXL inst_cellmath__24_0_I3598 (.Y(N8335), .A(N8328));
INVXL inst_cellmath__24_0_I3597 (.Y(N8334), .A(N8328));
XOR2XL inst_cellmath__24_0_I590 (.Y(N3033), .A(b_man[9]), .B(b_man[7]));
NAND2X2 inst_cellmath__24_0_I591 (.Y(N3114), .A(N3033), .B(N2779));
INVX1 inst_cellmath__24_0_I592 (.Y(N3564), .A(b_man[9]));
NAND2XL inst_cellmath__24_0_I593 (.Y(N2916), .A(b_man[7]), .B(b_man[8]));
AND2XL inst_cellmath__24_0_I594 (.Y(N3251), .A(b_man[9]), .B(N2916));
XNOR2X1 inst_cellmath__24_0_I595 (.Y(N2375), .A(N3445), .B(N3564));
OAI22XL inst_cellmath__24_0_I596 (.Y(N3586), .A0(N2375), .A1(N8335), .B0(N3564), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I597 (.Y(N3053), .A(N2228), .B(N3564));
OAI22XL inst_cellmath__24_0_I598 (.Y(N2718), .A0(N3053), .A1(N8335), .B0(N2375), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I599 (.Y(N2179), .A(N2573), .B(N3564));
OAI22XL inst_cellmath__24_0_I600 (.Y(N3400), .A0(N2179), .A1(N8334), .B0(N3053), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I601 (.Y(N2861), .A(N2911), .B(N3564));
OAI22XL inst_cellmath__24_0_I602 (.Y(N2520), .A0(N2861), .A1(N8334), .B0(N2179), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I603 (.Y(N3524), .A(N3243), .B(N3564));
OAI22XL inst_cellmath__24_0_I604 (.Y(N3193), .A0(N3524), .A1(N8334), .B0(N2861), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I605 (.Y(N2662), .A(N3578), .B(N3564));
OAI22XL inst_cellmath__24_0_I606 (.Y(N2318), .A0(N2662), .A1(N8334), .B0(N3524), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I607 (.Y(N3339), .A(N2368), .B(N3564));
OAI22XL inst_cellmath__24_0_I608 (.Y(N2996), .A0(N3339), .A1(N8334), .B0(N2662), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I609 (.Y(N2460), .A(N2713), .B(N3564));
OAI22XL inst_cellmath__24_0_I610 (.Y(N3667), .A0(N2460), .A1(N8334), .B0(N3339), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I611 (.Y(N3141), .A(N3047), .B(N3564));
OAI22XL inst_cellmath__24_0_I612 (.Y(N2806), .A0(N3141), .A1(N8334), .B0(N2460), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I613 (.Y(N2261), .A(N3391), .B(N3564));
OAI22XL inst_cellmath__24_0_I614 (.Y(N3470), .A0(N2261), .A1(N8334), .B0(N3141), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I615 (.Y(N2942), .A(N2171), .B(N3564));
OAI22XL inst_cellmath__24_0_I616 (.Y(N2603), .A0(N2942), .A1(N8335), .B0(N2261), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I617 (.Y(N3613), .A(N2511), .B(N3564));
OAI22XL inst_cellmath__24_0_I618 (.Y(N3278), .A0(N3613), .A1(N8335), .B0(N2942), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I619 (.Y(N2745), .A(N2853), .B(N3564));
OAI22XL inst_cellmath__24_0_I620 (.Y(N2399), .A0(N2745), .A1(N8335), .B0(N3613), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I621 (.Y(N3422), .A(N3186), .B(N3564));
OAI22XL inst_cellmath__24_0_I622 (.Y(N3080), .A0(N3422), .A1(N8335), .B0(N2745), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I623 (.Y(N2546), .A(N3513), .B(N3564));
OAI22XL inst_cellmath__24_0_I624 (.Y(N2201), .A0(N2546), .A1(N8334), .B0(N3422), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I625 (.Y(N3219), .A(N2308), .B(N3564));
OAI22XL inst_cellmath__24_0_I626 (.Y(N2886), .A0(N3219), .A1(N8334), .B0(N2546), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I627 (.Y(N2348), .A(N2653), .B(N3564));
OAI22XL inst_cellmath__24_0_I628 (.Y(N3551), .A0(N2348), .A1(N8334), .B0(N3219), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I629 (.Y(N3023), .A(N2987), .B(N3564));
OAI22XL inst_cellmath__24_0_I630 (.Y(N2688), .A0(N3023), .A1(N8334), .B0(N2348), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I631 (.Y(N2148), .A(N3329), .B(N3564));
OAI22XL inst_cellmath__24_0_I632 (.Y(N3363), .A0(N2148), .A1(N8334), .B0(N3023), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I633 (.Y(N2833), .A(N3660), .B(N3564));
OAI22XL inst_cellmath__24_0_I634 (.Y(N2484), .A0(N2833), .A1(N8334), .B0(N2148), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I635 (.Y(N3495), .A(N2452), .B(N3564));
OAI22XL inst_cellmath__24_0_I636 (.Y(N3166), .A0(N3495), .A1(N8334), .B0(N2833), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I637 (.Y(N2629), .A(N2799), .B(N3564));
OAI22XL inst_cellmath__24_0_I638 (.Y(N2287), .A0(N2629), .A1(N8334), .B0(N3495), .B1(N3114));
XNOR2X1 inst_cellmath__24_0_I639 (.Y(N3303), .A(N3134), .B(N3564));
OAI22XL inst_cellmath__24_0_I640 (.Y(N2967), .A0(N3303), .A1(N8335), .B0(N2629), .B1(N3114));
INVXL inst_cellmath__24_0_I641 (.Y(N2428), .A(N3564));
OAI22XL inst_cellmath__24_0_I642 (.Y(N3639), .A0(N2428), .A1(N8335), .B0(N3303), .B1(N3114));
MXI2XL inst_cellmath__24_0_I643 (.Y(N2772), .A(N3114), .B(N8335), .S0(N2428));
XNOR2X1 inst_cellmath__24_0_I644 (.Y(N2712), .A(b_man[10]), .B(b_man[9]));
INVXL inst_cellmath__24_0_I3599 (.Y(N8336), .A(N2712));
INVXL inst_cellmath__24_0_I3606 (.Y(N8343), .A(N8336));
INVXL inst_cellmath__24_0_I3605 (.Y(N8342), .A(N8336));
XOR2XL inst_cellmath__24_0_I645 (.Y(N2267), .A(b_man[11]), .B(b_man[9]));
NAND2X2 inst_cellmath__24_0_I646 (.Y(N3048), .A(N2267), .B(N2712));
INVX1 inst_cellmath__24_0_I647 (.Y(N3258), .A(b_man[11]));
NAND2XL inst_cellmath__24_0_I648 (.Y(N2855), .A(b_man[9]), .B(b_man[10]));
AND2XL inst_cellmath__24_0_I649 (.Y(N3185), .A(b_man[11]), .B(N2855));
XNOR2X1 inst_cellmath__24_0_I650 (.Y(N2311), .A(N3445), .B(N3258));
OAI22XL inst_cellmath__24_0_I651 (.Y(N3515), .A0(N2311), .A1(N8343), .B0(N3258), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I652 (.Y(N2989), .A(N2228), .B(N3258));
OAI22XL inst_cellmath__24_0_I653 (.Y(N2652), .A0(N2989), .A1(N8343), .B0(N2311), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I654 (.Y(N3659), .A(N2573), .B(N3258));
OAI22XL inst_cellmath__24_0_I655 (.Y(N3331), .A0(N3659), .A1(N8342), .B0(N2989), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I656 (.Y(N2800), .A(N2911), .B(N3258));
OAI22XL inst_cellmath__24_0_I657 (.Y(N2453), .A0(N2800), .A1(N8342), .B0(N3659), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I658 (.Y(N3465), .A(N3243), .B(N3258));
OAI22XL inst_cellmath__24_0_I659 (.Y(N3133), .A0(N3465), .A1(N8342), .B0(N2800), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I660 (.Y(N2596), .A(N3578), .B(N3258));
OAI22XL inst_cellmath__24_0_I661 (.Y(N2255), .A0(N2596), .A1(N8342), .B0(N3465), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I662 (.Y(N3273), .A(N2368), .B(N3258));
OAI22XL inst_cellmath__24_0_I663 (.Y(N2937), .A0(N3273), .A1(N8343), .B0(N2596), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I664 (.Y(N2393), .A(N2713), .B(N3258));
OAI22XL inst_cellmath__24_0_I665 (.Y(N3607), .A0(N2393), .A1(N8343), .B0(N3273), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I666 (.Y(N3072), .A(N3047), .B(N3258));
OAI22XL inst_cellmath__24_0_I667 (.Y(N2738), .A0(N3072), .A1(N8343), .B0(N2393), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I668 (.Y(N2194), .A(N3391), .B(N3258));
OAI22XL inst_cellmath__24_0_I669 (.Y(N3416), .A0(N2194), .A1(N8343), .B0(N3072), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I670 (.Y(N2879), .A(N2171), .B(N3258));
OAI22XL inst_cellmath__24_0_I671 (.Y(N2539), .A0(N2879), .A1(N8343), .B0(N2194), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I672 (.Y(N3542), .A(N2511), .B(N3258));
OAI22XL inst_cellmath__24_0_I673 (.Y(N3213), .A0(N3542), .A1(N8343), .B0(N2879), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I674 (.Y(N2683), .A(N2853), .B(N3258));
OAI22XL inst_cellmath__24_0_I675 (.Y(N2341), .A0(N2683), .A1(N8343), .B0(N3542), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I676 (.Y(N3358), .A(N3186), .B(N3258));
OAI22XL inst_cellmath__24_0_I677 (.Y(N3016), .A0(N3358), .A1(N8343), .B0(N2683), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I678 (.Y(N2476), .A(N3513), .B(N3258));
OAI22XL inst_cellmath__24_0_I679 (.Y(N3686), .A0(N2476), .A1(N8342), .B0(N3358), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I680 (.Y(N3160), .A(N2308), .B(N3258));
OAI22XL inst_cellmath__24_0_I681 (.Y(N2822), .A0(N3160), .A1(N8342), .B0(N2476), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I682 (.Y(N2279), .A(N2653), .B(N3258));
OAI22XL inst_cellmath__24_0_I683 (.Y(N3485), .A0(N2279), .A1(N8342), .B0(N3160), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I684 (.Y(N2957), .A(N2987), .B(N3258));
OAI22XL inst_cellmath__24_0_I685 (.Y(N2623), .A0(N2957), .A1(N8342), .B0(N2279), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I686 (.Y(N3633), .A(N3329), .B(N3258));
OAI22XL inst_cellmath__24_0_I687 (.Y(N3297), .A0(N3633), .A1(N8342), .B0(N2957), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I688 (.Y(N2765), .A(N3660), .B(N3258));
OAI22XL inst_cellmath__24_0_I689 (.Y(N2418), .A0(N2765), .A1(N8342), .B0(N3633), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I690 (.Y(N3439), .A(N2452), .B(N3258));
OAI22XL inst_cellmath__24_0_I691 (.Y(N3103), .A0(N3439), .A1(N8342), .B0(N2765), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I692 (.Y(N2567), .A(N2799), .B(N3258));
OAI22XL inst_cellmath__24_0_I693 (.Y(N2222), .A0(N2567), .A1(N8342), .B0(N3439), .B1(N3048));
XNOR2X1 inst_cellmath__24_0_I694 (.Y(N3237), .A(N3134), .B(N3258));
OAI22XL inst_cellmath__24_0_I695 (.Y(N2903), .A0(N3237), .A1(N8342), .B0(N2567), .B1(N3048));
INVXL inst_cellmath__24_0_I696 (.Y(N2364), .A(N3258));
OAI22XL inst_cellmath__24_0_I697 (.Y(N3573), .A0(N2364), .A1(N8342), .B0(N3237), .B1(N3048));
MXI2XL inst_cellmath__24_0_I698 (.Y(N2706), .A(N3048), .B(N8342), .S0(N2364));
XNOR2X1 inst_cellmath__24_0_I699 (.Y(N2646), .A(b_man[12]), .B(b_man[11]));
XOR2XL inst_cellmath__24_0_I700 (.Y(N3060), .A(b_man[13]), .B(b_man[11]));
NAND2X2 inst_cellmath__24_0_I701 (.Y(N2981), .A(N3060), .B(N2646));
INVX1 inst_cellmath__24_0_I702 (.Y(N2947), .A(b_man[13]));
NAND2XL inst_cellmath__24_0_I703 (.Y(N2795), .A(b_man[11]), .B(b_man[12]));
AND2XL inst_cellmath__24_0_I704 (.Y(N3126), .A(b_man[13]), .B(N2795));
XNOR2X1 inst_cellmath__24_0_I705 (.Y(N2248), .A(N3445), .B(N2947));
OAI22XL inst_cellmath__24_0_I706 (.Y(N3460), .A0(N2248), .A1(N2646), .B0(N2947), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I707 (.Y(N2929), .A(N2228), .B(N2947));
OAI22XL inst_cellmath__24_0_I708 (.Y(N2592), .A0(N2929), .A1(N2646), .B0(N2248), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I709 (.Y(N3597), .A(N2573), .B(N2947));
OAI22XL inst_cellmath__24_0_I710 (.Y(N3267), .A0(N3597), .A1(N2646), .B0(N2929), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I711 (.Y(N2731), .A(N2911), .B(N2947));
OAI22XL inst_cellmath__24_0_I712 (.Y(N2387), .A0(N2731), .A1(N2646), .B0(N3597), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I713 (.Y(N3410), .A(N3243), .B(N2947));
OAI22XL inst_cellmath__24_0_I714 (.Y(N3065), .A0(N3410), .A1(N2646), .B0(N2731), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I715 (.Y(N2533), .A(N3578), .B(N2947));
OAI22XL inst_cellmath__24_0_I716 (.Y(N2189), .A0(N2533), .A1(N2646), .B0(N3410), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I717 (.Y(N3206), .A(N2368), .B(N2947));
OAI22XL inst_cellmath__24_0_I718 (.Y(N2873), .A0(N3206), .A1(N2646), .B0(N2533), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I719 (.Y(N2334), .A(N2713), .B(N2947));
OAI22XL inst_cellmath__24_0_I720 (.Y(N3535), .A0(N2334), .A1(N2646), .B0(N3206), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I721 (.Y(N3008), .A(N3047), .B(N2947));
OAI22XL inst_cellmath__24_0_I722 (.Y(N2675), .A0(N3008), .A1(N2646), .B0(N2334), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I723 (.Y(N3678), .A(N3391), .B(N2947));
OAI22XL inst_cellmath__24_0_I724 (.Y(N3348), .A0(N3678), .A1(N2646), .B0(N3008), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I725 (.Y(N2816), .A(N2171), .B(N2947));
OAI22XL inst_cellmath__24_0_I726 (.Y(N2470), .A0(N2816), .A1(N2646), .B0(N3678), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I727 (.Y(N3478), .A(N2511), .B(N2947));
OAI22XL inst_cellmath__24_0_I728 (.Y(N3151), .A0(N3478), .A1(N2646), .B0(N2816), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I729 (.Y(N2613), .A(N2853), .B(N2947));
OAI22XL inst_cellmath__24_0_I730 (.Y(N2272), .A0(N2613), .A1(N2646), .B0(N3478), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I731 (.Y(N3289), .A(N3186), .B(N2947));
OAI22XL inst_cellmath__24_0_I732 (.Y(N2952), .A0(N3289), .A1(N2646), .B0(N2613), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I733 (.Y(N2410), .A(N3513), .B(N2947));
OAI22XL inst_cellmath__24_0_I734 (.Y(N3625), .A0(N2410), .A1(N2646), .B0(N3289), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I735 (.Y(N3094), .A(N2308), .B(N2947));
OAI22XL inst_cellmath__24_0_I736 (.Y(N2758), .A0(N3094), .A1(N2646), .B0(N2410), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I737 (.Y(N2214), .A(N2653), .B(N2947));
OAI22XL inst_cellmath__24_0_I738 (.Y(N3432), .A0(N2214), .A1(N2646), .B0(N3094), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I739 (.Y(N2894), .A(N2987), .B(N2947));
OAI22XL inst_cellmath__24_0_I740 (.Y(N2559), .A0(N2894), .A1(N2646), .B0(N2214), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I741 (.Y(N3567), .A(N3329), .B(N2947));
OAI22XL inst_cellmath__24_0_I742 (.Y(N3229), .A0(N3567), .A1(N2646), .B0(N2894), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I743 (.Y(N2699), .A(N3660), .B(N2947));
OAI22XL inst_cellmath__24_0_I744 (.Y(N2359), .A0(N2699), .A1(N2646), .B0(N3567), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I745 (.Y(N3373), .A(N2452), .B(N2947));
OAI22XL inst_cellmath__24_0_I746 (.Y(N3035), .A0(N3373), .A1(N2646), .B0(N2699), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I747 (.Y(N2497), .A(N2799), .B(N2947));
OAI22XL inst_cellmath__24_0_I748 (.Y(N2159), .A0(N2497), .A1(N2646), .B0(N3373), .B1(N2981));
XNOR2X1 inst_cellmath__24_0_I749 (.Y(N3173), .A(N3134), .B(N2947));
OAI22XL inst_cellmath__24_0_I750 (.Y(N2843), .A0(N3173), .A1(N2646), .B0(N2497), .B1(N2981));
INVXL inst_cellmath__24_0_I751 (.Y(N2296), .A(N2947));
OAI22XL inst_cellmath__24_0_I752 (.Y(N3504), .A0(N2296), .A1(N2646), .B0(N3173), .B1(N2981));
MXI2XL inst_cellmath__24_0_I753 (.Y(N2639), .A(N2981), .B(N2646), .S0(N2296));
XNOR2X1 inst_cellmath__24_0_I754 (.Y(N2586), .A(b_man[14]), .B(b_man[13]));
INVXL inst_cellmath__24_0_I3615 (.Y(N8352), .A(N2586));
INVXL inst_cellmath__24_0_I3622 (.Y(N8359), .A(N8352));
INVXL inst_cellmath__24_0_I3621 (.Y(N8358), .A(N8352));
XOR2XL inst_cellmath__24_0_I755 (.Y(N2295), .A(b_man[15]), .B(b_man[13]));
NAND2X1 inst_cellmath__24_0_I756 (.Y(N2923), .A(N2295), .B(N2586));
INVX1 inst_cellmath__24_0_I757 (.Y(N2352), .A(b_man[15]));
NAND2XL inst_cellmath__24_0_I758 (.Y(N2721), .A(b_man[13]), .B(b_man[14]));
AND2XL inst_cellmath__24_0_I759 (.Y(N3058), .A(b_man[15]), .B(N2721));
XNOR2X1 inst_cellmath__24_0_I760 (.Y(N2184), .A(N3445), .B(N2352));
OAI22XL inst_cellmath__24_0_I761 (.Y(N3403), .A0(N2184), .A1(N8359), .B0(N2352), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I762 (.Y(N2865), .A(N2228), .B(N2352));
OAI22XL inst_cellmath__24_0_I763 (.Y(N2523), .A0(N2865), .A1(N8359), .B0(N2184), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I764 (.Y(N3528), .A(N2573), .B(N2352));
OAI22XL inst_cellmath__24_0_I765 (.Y(N3200), .A0(N3528), .A1(N8358), .B0(N2865), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I766 (.Y(N2667), .A(N2911), .B(N2352));
OAI22XL inst_cellmath__24_0_I767 (.Y(N2323), .A0(N2667), .A1(N8358), .B0(N3528), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I768 (.Y(N3342), .A(N3243), .B(N2352));
OAI22XL inst_cellmath__24_0_I769 (.Y(N2999), .A0(N3342), .A1(N8358), .B0(N2667), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I770 (.Y(N2463), .A(N3578), .B(N2352));
OAI22XL inst_cellmath__24_0_I771 (.Y(N3672), .A0(N2463), .A1(N8358), .B0(N3342), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I772 (.Y(N3146), .A(N2368), .B(N2352));
OAI22XL inst_cellmath__24_0_I773 (.Y(N2811), .A0(N3146), .A1(N8359), .B0(N2463), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I774 (.Y(N2264), .A(N2713), .B(N2352));
OAI22XL inst_cellmath__24_0_I775 (.Y(N3472), .A0(N2264), .A1(N8359), .B0(N3146), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I776 (.Y(N2946), .A(N3047), .B(N2352));
OAI22XL inst_cellmath__24_0_I777 (.Y(N2606), .A0(N2946), .A1(N8359), .B0(N2264), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I778 (.Y(N3618), .A(N3391), .B(N2352));
OAI22XL inst_cellmath__24_0_I779 (.Y(N3282), .A0(N3618), .A1(N8359), .B0(N2946), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I780 (.Y(N2751), .A(N2171), .B(N2352));
OAI22XL inst_cellmath__24_0_I781 (.Y(N2403), .A0(N2751), .A1(N8358), .B0(N3618), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I782 (.Y(N3426), .A(N2511), .B(N2352));
OAI22XL inst_cellmath__24_0_I783 (.Y(N3087), .A0(N3426), .A1(N8358), .B0(N2751), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I784 (.Y(N2554), .A(N2853), .B(N2352));
OAI22XL inst_cellmath__24_0_I785 (.Y(N2206), .A0(N2554), .A1(N8358), .B0(N3426), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I786 (.Y(N3223), .A(N3186), .B(N2352));
OAI22XL inst_cellmath__24_0_I787 (.Y(N2890), .A0(N3223), .A1(N8358), .B0(N2554), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I788 (.Y(N2351), .A(N3513), .B(N2352));
OAI22XL inst_cellmath__24_0_I789 (.Y(N3556), .A0(N2351), .A1(N8359), .B0(N3223), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I790 (.Y(N3028), .A(N2308), .B(N2352));
OAI22XL inst_cellmath__24_0_I791 (.Y(N2693), .A0(N3028), .A1(N8359), .B0(N2351), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I792 (.Y(N2153), .A(N2653), .B(N2352));
OAI22XL inst_cellmath__24_0_I793 (.Y(N3366), .A0(N2153), .A1(N8359), .B0(N3028), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I794 (.Y(N2836), .A(N2987), .B(N2352));
OAI22XL inst_cellmath__24_0_I795 (.Y(N2490), .A0(N2836), .A1(N8359), .B0(N2153), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I796 (.Y(N3498), .A(N3329), .B(N2352));
OAI22XL inst_cellmath__24_0_I797 (.Y(N3168), .A0(N3498), .A1(N8359), .B0(N2836), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I798 (.Y(N2634), .A(N3660), .B(N2352));
OAI22XL inst_cellmath__24_0_I799 (.Y(N2291), .A0(N2634), .A1(N8359), .B0(N3498), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I800 (.Y(N3307), .A(N2452), .B(N2352));
OAI22XL inst_cellmath__24_0_I801 (.Y(N2972), .A0(N3307), .A1(N8359), .B0(N2634), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I802 (.Y(N2432), .A(N2799), .B(N2352));
OAI22XL inst_cellmath__24_0_I803 (.Y(N3643), .A0(N2432), .A1(N8359), .B0(N3307), .B1(N2923));
XNOR2X1 inst_cellmath__24_0_I804 (.Y(N3112), .A(N3134), .B(N2352));
OAI22XL inst_cellmath__24_0_I805 (.Y(N2775), .A0(N3112), .A1(N8358), .B0(N2432), .B1(N2923));
INVXL inst_cellmath__24_0_I806 (.Y(N2232), .A(N2352));
OAI22XL inst_cellmath__24_0_I807 (.Y(N3449), .A0(N2232), .A1(N8358), .B0(N3112), .B1(N2923));
MXI2XL inst_cellmath__24_0_I808 (.Y(N2580), .A(N2923), .B(N8358), .S0(N2232));
XNOR2X1 inst_cellmath__24_0_I809 (.Y(N2519), .A(b_man[16]), .B(b_man[15]));
XOR2XL inst_cellmath__24_0_I810 (.Y(N3090), .A(b_man[17]), .B(b_man[15]));
NAND2X2 inst_cellmath__24_0_I811 (.Y(N2860), .A(N3090), .B(N2519));
INVX1 inst_cellmath__24_0_I812 (.Y(N3583), .A(b_man[17]));
NAND2XL inst_cellmath__24_0_I813 (.Y(N2658), .A(b_man[15]), .B(b_man[16]));
AND2XL inst_cellmath__24_0_I814 (.Y(N2994), .A(b_man[17]), .B(N2658));
XNOR2X1 inst_cellmath__24_0_I815 (.Y(N3665), .A(N3445), .B(N3583));
OAI22XL inst_cellmath__24_0_I816 (.Y(N3336), .A0(N3665), .A1(N2519), .B0(N3583), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I817 (.Y(N2804), .A(N2228), .B(N3583));
OAI22XL inst_cellmath__24_0_I818 (.Y(N2458), .A0(N2804), .A1(N2519), .B0(N3665), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I819 (.Y(N3468), .A(N2573), .B(N3583));
OAI22XL inst_cellmath__24_0_I820 (.Y(N3137), .A0(N3468), .A1(N2519), .B0(N2804), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I821 (.Y(N2600), .A(N2911), .B(N3583));
OAI22XL inst_cellmath__24_0_I822 (.Y(N2259), .A0(N2600), .A1(N2519), .B0(N3468), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I823 (.Y(N3276), .A(N3243), .B(N3583));
OAI22XL inst_cellmath__24_0_I824 (.Y(N2941), .A0(N3276), .A1(N2519), .B0(N2600), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I825 (.Y(N2397), .A(N3578), .B(N3583));
OAI22XL inst_cellmath__24_0_I826 (.Y(N3612), .A0(N2397), .A1(N2519), .B0(N3276), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I827 (.Y(N3079), .A(N2368), .B(N3583));
OAI22XL inst_cellmath__24_0_I828 (.Y(N2743), .A0(N3079), .A1(N2519), .B0(N2397), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I829 (.Y(N2199), .A(N2713), .B(N3583));
OAI22XL inst_cellmath__24_0_I830 (.Y(N3419), .A0(N2199), .A1(N2519), .B0(N3079), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I831 (.Y(N2882), .A(N3047), .B(N3583));
OAI22XL inst_cellmath__24_0_I832 (.Y(N2545), .A0(N2882), .A1(N2519), .B0(N2199), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I833 (.Y(N3550), .A(N3391), .B(N3583));
OAI22XL inst_cellmath__24_0_I834 (.Y(N3217), .A0(N3550), .A1(N2519), .B0(N2882), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I835 (.Y(N2686), .A(N2171), .B(N3583));
OAI22XL inst_cellmath__24_0_I836 (.Y(N2345), .A0(N2686), .A1(N2519), .B0(N3550), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I837 (.Y(N3362), .A(N2511), .B(N3583));
OAI22XL inst_cellmath__24_0_I838 (.Y(N3021), .A0(N3362), .A1(N2519), .B0(N2686), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I839 (.Y(N2483), .A(N2853), .B(N3583));
OAI22XL inst_cellmath__24_0_I840 (.Y(N3689), .A0(N2483), .A1(N2519), .B0(N3362), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I841 (.Y(N3164), .A(N3186), .B(N3583));
OAI22XL inst_cellmath__24_0_I842 (.Y(N2829), .A0(N3164), .A1(N2519), .B0(N2483), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I843 (.Y(N2284), .A(N3513), .B(N3583));
OAI22XL inst_cellmath__24_0_I844 (.Y(N3492), .A0(N2284), .A1(N2519), .B0(N3164), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I845 (.Y(N2965), .A(N2308), .B(N3583));
OAI22XL inst_cellmath__24_0_I846 (.Y(N2626), .A0(N2965), .A1(N2519), .B0(N2284), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I847 (.Y(N3637), .A(N2653), .B(N3583));
OAI22XL inst_cellmath__24_0_I848 (.Y(N3300), .A0(N3637), .A1(N2519), .B0(N2965), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I849 (.Y(N2768), .A(N2987), .B(N3583));
OAI22XL inst_cellmath__24_0_I850 (.Y(N2425), .A0(N2768), .A1(N2519), .B0(N3637), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I851 (.Y(N3444), .A(N3329), .B(N3583));
OAI22XL inst_cellmath__24_0_I852 (.Y(N3107), .A0(N3444), .A1(N2519), .B0(N2768), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I853 (.Y(N2572), .A(N3660), .B(N3583));
OAI22XL inst_cellmath__24_0_I854 (.Y(N2225), .A0(N2572), .A1(N2519), .B0(N3444), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I855 (.Y(N3240), .A(N2452), .B(N3583));
OAI22XL inst_cellmath__24_0_I856 (.Y(N2910), .A0(N3240), .A1(N2519), .B0(N2572), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I857 (.Y(N2367), .A(N2799), .B(N3583));
OAI22XL inst_cellmath__24_0_I858 (.Y(N3576), .A0(N2367), .A1(N2519), .B0(N3240), .B1(N2860));
XNOR2X1 inst_cellmath__24_0_I859 (.Y(N3046), .A(N3134), .B(N3583));
OAI22XL inst_cellmath__24_0_I860 (.Y(N2710), .A0(N3046), .A1(N2519), .B0(N2367), .B1(N2860));
INVXL inst_cellmath__24_0_I861 (.Y(N2169), .A(N3583));
OAI22XL inst_cellmath__24_0_I862 (.Y(N3390), .A0(N2169), .A1(N2519), .B0(N3046), .B1(N2860));
MXI2XL inst_cellmath__24_0_I863 (.Y(N2509), .A(N2860), .B(N2519), .S0(N2169));
XNOR2X1 inst_cellmath__24_0_I864 (.Y(N2450), .A(b_man[18]), .B(b_man[17]));
XOR2XL inst_cellmath__24_0_I865 (.Y(N2325), .A(b_man[19]), .B(b_man[17]));
NAND2X1 inst_cellmath__24_0_I866 (.Y(N2659), .A(N2325), .B(N2450));
INVXL inst_cellmath__24_0_I867 (.Y(N2993), .A(b_man[19]));
NAND2XL inst_cellmath__24_0_I868 (.Y(N2595), .A(b_man[17]), .B(b_man[18]));
AND2XL inst_cellmath__24_0_I869 (.Y(N2933), .A(b_man[19]), .B(N2595));
XNOR2X1 inst_cellmath__24_0_I870 (.Y(N3603), .A(N3445), .B(N2993));
OAI22XL inst_cellmath__24_0_I871 (.Y(N3271), .A0(N3603), .A1(N2450), .B0(N2993), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I872 (.Y(N2736), .A(N2228), .B(N2993));
OAI22XL inst_cellmath__24_0_I873 (.Y(N2392), .A0(N2736), .A1(N2450), .B0(N3603), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I874 (.Y(N3413), .A(N2573), .B(N2993));
OAI22XL inst_cellmath__24_0_I875 (.Y(N3070), .A0(N3413), .A1(N2450), .B0(N2736), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I876 (.Y(N2537), .A(N2911), .B(N2993));
OAI22XL inst_cellmath__24_0_I877 (.Y(N2192), .A0(N2537), .A1(N2450), .B0(N3413), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I878 (.Y(N3211), .A(N3243), .B(N2993));
OAI22XL inst_cellmath__24_0_I879 (.Y(N2877), .A0(N3211), .A1(N2450), .B0(N2537), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I880 (.Y(N2338), .A(N3578), .B(N2993));
OAI22XL inst_cellmath__24_0_I881 (.Y(N3538), .A0(N2338), .A1(N2450), .B0(N3211), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I882 (.Y(N3013), .A(N2368), .B(N2993));
OAI22XL inst_cellmath__24_0_I883 (.Y(N2680), .A0(N3013), .A1(N2450), .B0(N2338), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I884 (.Y(N3684), .A(N2713), .B(N2993));
OAI22XL inst_cellmath__24_0_I885 (.Y(N3355), .A0(N3684), .A1(N2450), .B0(N3013), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I886 (.Y(N2820), .A(N3047), .B(N2993));
OAI22XL inst_cellmath__24_0_I887 (.Y(N2474), .A0(N2820), .A1(N2450), .B0(N3684), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I888 (.Y(N3482), .A(N3391), .B(N2993));
OAI22XL inst_cellmath__24_0_I889 (.Y(N3156), .A0(N3482), .A1(N2450), .B0(N2820), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I890 (.Y(N2618), .A(N2171), .B(N2993));
OAI22XL inst_cellmath__24_0_I891 (.Y(N2277), .A0(N2618), .A1(N2450), .B0(N3482), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I892 (.Y(N3292), .A(N2511), .B(N2993));
OAI22XL inst_cellmath__24_0_I893 (.Y(N2956), .A0(N3292), .A1(N2450), .B0(N2618), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I894 (.Y(N2417), .A(N2853), .B(N2993));
OAI22XL inst_cellmath__24_0_I895 (.Y(N3630), .A0(N2417), .A1(N2450), .B0(N3292), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I896 (.Y(N3099), .A(N3186), .B(N2993));
OAI22XL inst_cellmath__24_0_I897 (.Y(N2762), .A0(N3099), .A1(N2450), .B0(N2417), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I898 (.Y(N2218), .A(N3513), .B(N2993));
OAI22XL inst_cellmath__24_0_I899 (.Y(N3438), .A0(N2218), .A1(N2450), .B0(N3099), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I900 (.Y(N2902), .A(N2308), .B(N2993));
OAI22XL inst_cellmath__24_0_I901 (.Y(N2564), .A0(N2902), .A1(N2450), .B0(N2218), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I902 (.Y(N3570), .A(N2653), .B(N2993));
OAI22XL inst_cellmath__24_0_I903 (.Y(N3234), .A0(N3570), .A1(N2450), .B0(N2902), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I904 (.Y(N2703), .A(N2987), .B(N2993));
OAI22XL inst_cellmath__24_0_I905 (.Y(N2363), .A0(N2703), .A1(N2450), .B0(N3570), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I906 (.Y(N3381), .A(N3329), .B(N2993));
OAI22XL inst_cellmath__24_0_I907 (.Y(N3039), .A0(N3381), .A1(N2450), .B0(N2703), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I908 (.Y(N2502), .A(N3660), .B(N2993));
OAI22XL inst_cellmath__24_0_I909 (.Y(N2163), .A0(N2502), .A1(N2450), .B0(N3381), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I910 (.Y(N3177), .A(N2452), .B(N2993));
OAI22XL inst_cellmath__24_0_I911 (.Y(N2847), .A0(N3177), .A1(N2450), .B0(N2502), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I912 (.Y(N2300), .A(N2799), .B(N2993));
OAI22XL inst_cellmath__24_0_I913 (.Y(N3507), .A0(N2300), .A1(N2450), .B0(N3177), .B1(N2659));
XNOR2X1 inst_cellmath__24_0_I914 (.Y(N2979), .A(N3134), .B(N2993));
OAI22XL inst_cellmath__24_0_I915 (.Y(N2642), .A0(N2979), .A1(N2450), .B0(N2300), .B1(N2659));
INVXL inst_cellmath__24_0_I916 (.Y(N3652), .A(N2993));
OAI22XL inst_cellmath__24_0_I917 (.Y(N3321), .A0(N3652), .A1(N2450), .B0(N2979), .B1(N2659));
MXI2XL inst_cellmath__24_0_I918 (.Y(N2442), .A(N2659), .B(N2450), .S0(N3652));
XNOR2X1 inst_cellmath__24_0_I919 (.Y(N2385), .A(b_man[20]), .B(b_man[19]));
XOR2XL inst_cellmath__24_0_I920 (.Y(N3118), .A(b_man[21]), .B(b_man[19]));
NAND2X1 inst_cellmath__24_0_I921 (.Y(N3609), .A(N3118), .B(N2385));
INVXL inst_cellmath__24_0_I922 (.Y(N2395), .A(b_man[21]));
NAND2XL inst_cellmath__24_0_I923 (.Y(N2529), .A(b_man[19]), .B(b_man[20]));
AND2XL inst_cellmath__24_0_I924 (.Y(N2871), .A(b_man[21]), .B(N2529));
XNOR2X1 inst_cellmath__24_0_I925 (.Y(N3533), .A(N3445), .B(N2395));
OAI22XL inst_cellmath__24_0_I926 (.Y(N3204), .A0(N3533), .A1(N2385), .B0(N2395), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I927 (.Y(N2673), .A(N2228), .B(N2395));
OAI22XL inst_cellmath__24_0_I928 (.Y(N2330), .A0(N2673), .A1(N2385), .B0(N3533), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I929 (.Y(N3346), .A(N2573), .B(N2395));
OAI22XL inst_cellmath__24_0_I930 (.Y(N3005), .A0(N3346), .A1(N2385), .B0(N2673), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I931 (.Y(N2468), .A(N2911), .B(N2395));
OAI22XL inst_cellmath__24_0_I932 (.Y(N3676), .A0(N2468), .A1(N2385), .B0(N3346), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I933 (.Y(N3150), .A(N3243), .B(N2395));
OAI22XL inst_cellmath__24_0_I934 (.Y(N2814), .A0(N3150), .A1(N2385), .B0(N2468), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I935 (.Y(N2270), .A(N3578), .B(N2395));
OAI22XL inst_cellmath__24_0_I936 (.Y(N3476), .A0(N2270), .A1(N2385), .B0(N3150), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I937 (.Y(N2950), .A(N2368), .B(N2395));
OAI22XL inst_cellmath__24_0_I938 (.Y(N2611), .A0(N2950), .A1(N2385), .B0(N2270), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I939 (.Y(N3622), .A(N2713), .B(N2395));
OAI22XL inst_cellmath__24_0_I940 (.Y(N3287), .A0(N3622), .A1(N2385), .B0(N2950), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I941 (.Y(N2757), .A(N3047), .B(N2395));
OAI22XL inst_cellmath__24_0_I942 (.Y(N2408), .A0(N2757), .A1(N2385), .B0(N3622), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I943 (.Y(N3430), .A(N3391), .B(N2395));
OAI22XL inst_cellmath__24_0_I944 (.Y(N3093), .A0(N3430), .A1(N2385), .B0(N2757), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I945 (.Y(N2557), .A(N2171), .B(N2395));
OAI22XL inst_cellmath__24_0_I946 (.Y(N2210), .A0(N2557), .A1(N2385), .B0(N3430), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I947 (.Y(N3227), .A(N2511), .B(N2395));
OAI22XL inst_cellmath__24_0_I948 (.Y(N2893), .A0(N3227), .A1(N2385), .B0(N2557), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I949 (.Y(N2356), .A(N2853), .B(N2395));
OAI22XL inst_cellmath__24_0_I950 (.Y(N3562), .A0(N2356), .A1(N2385), .B0(N3227), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I951 (.Y(N3032), .A(N3186), .B(N2395));
OAI22XL inst_cellmath__24_0_I952 (.Y(N2697), .A0(N3032), .A1(N2385), .B0(N2356), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I953 (.Y(N2157), .A(N3513), .B(N2395));
OAI22XL inst_cellmath__24_0_I954 (.Y(N3371), .A0(N2157), .A1(N2385), .B0(N3032), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I955 (.Y(N2841), .A(N2308), .B(N2395));
OAI22XL inst_cellmath__24_0_I956 (.Y(N2495), .A0(N2841), .A1(N2385), .B0(N2157), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I957 (.Y(N3502), .A(N2653), .B(N2395));
OAI22XL inst_cellmath__24_0_I958 (.Y(N3172), .A0(N3502), .A1(N2385), .B0(N2841), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I959 (.Y(N2635), .A(N2987), .B(N2395));
OAI22XL inst_cellmath__24_0_I960 (.Y(N2294), .A0(N2635), .A1(N2385), .B0(N3502), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I961 (.Y(N3314), .A(N3329), .B(N2395));
OAI22XL inst_cellmath__24_0_I962 (.Y(N2974), .A0(N3314), .A1(N2385), .B0(N2635), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I963 (.Y(N2436), .A(N3660), .B(N2395));
OAI22XL inst_cellmath__24_0_I964 (.Y(N3646), .A0(N2436), .A1(N2385), .B0(N3314), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I965 (.Y(N3115), .A(N2452), .B(N2395));
OAI22XL inst_cellmath__24_0_I966 (.Y(N2783), .A0(N3115), .A1(N2385), .B0(N2436), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I967 (.Y(N2238), .A(N2799), .B(N2395));
OAI22XL inst_cellmath__24_0_I968 (.Y(N3451), .A0(N2238), .A1(N2385), .B0(N3115), .B1(N3609));
XNOR2X1 inst_cellmath__24_0_I969 (.Y(N2919), .A(N3134), .B(N2395));
OAI22XL inst_cellmath__24_0_I970 (.Y(N2583), .A0(N2919), .A1(N2385), .B0(N2238), .B1(N3609));
INVXL inst_cellmath__24_0_I971 (.Y(N3587), .A(N2395));
OAI22XL inst_cellmath__24_0_I972 (.Y(N3256), .A0(N3587), .A1(N2385), .B0(N2919), .B1(N3609));
MXI2XL inst_cellmath__24_0_I973 (.Y(N2377), .A(N3609), .B(N2385), .S0(N3587));
XNOR2X1 inst_cellmath__24_0_I974 (.Y(N2320), .A(b_man[22]), .B(b_man[21]));
OR2XL inst_cellmath__24_0_I975 (.Y(N2963), .A(b_man[22]), .B(b_man[21]));
NAND2XL inst_cellmath__24_0_I976 (.Y(N2807), .A(b_man[21]), .B(b_man[22]));
INVXL inst_cellmath__24_0_I977 (.Y(N2748), .A(N3445));
OAI21XL inst_cellmath__24_0_I978 (.Y(N2400), .A0(N2320), .A1(N2748), .B0(N2963));
INVXL inst_cellmath__24_0_I979 (.Y(N3423), .A(N2228));
OAI22XL inst_cellmath__24_0_I980 (.Y(N3085), .A0(N3423), .A1(N2320), .B0(N2748), .B1(N2963));
INVXL inst_cellmath__24_0_I981 (.Y(N2550), .A(N2573));
OAI22XL inst_cellmath__24_0_I982 (.Y(N2203), .A0(N2550), .A1(N2320), .B0(N3423), .B1(N2963));
INVXL inst_cellmath__24_0_I983 (.Y(N3220), .A(N2911));
OAI22XL inst_cellmath__24_0_I984 (.Y(N2887), .A0(N3220), .A1(N2320), .B0(N2550), .B1(N2963));
INVXL inst_cellmath__24_0_I985 (.Y(N2349), .A(N3243));
OAI22XL inst_cellmath__24_0_I986 (.Y(N3554), .A0(N2349), .A1(N2320), .B0(N3220), .B1(N2963));
INVXL inst_cellmath__24_0_I987 (.Y(N3026), .A(N3578));
OAI22XL inst_cellmath__24_0_I988 (.Y(N2690), .A0(N3026), .A1(N2320), .B0(N2349), .B1(N2963));
INVXL inst_cellmath__24_0_I989 (.Y(N2150), .A(N2368));
OAI22XL inst_cellmath__24_0_I990 (.Y(N3364), .A0(N2150), .A1(N2320), .B0(N3026), .B1(N2963));
INVXL inst_cellmath__24_0_I991 (.Y(N2835), .A(N2713));
OAI22XL inst_cellmath__24_0_I992 (.Y(N2487), .A0(N2835), .A1(N2320), .B0(N2150), .B1(N2963));
INVXL inst_cellmath__24_0_I993 (.Y(N3497), .A(N3047));
OAI22XL inst_cellmath__24_0_I994 (.Y(N3167), .A0(N3497), .A1(N2320), .B0(N2835), .B1(N2963));
INVXL inst_cellmath__24_0_I995 (.Y(N2631), .A(N3391));
OAI22XL inst_cellmath__24_0_I996 (.Y(N2288), .A0(N2631), .A1(N2320), .B0(N3497), .B1(N2963));
INVXL inst_cellmath__24_0_I997 (.Y(N3305), .A(N2171));
OAI22XL inst_cellmath__24_0_I998 (.Y(N2970), .A0(N3305), .A1(N2320), .B0(N2631), .B1(N2963));
INVXL inst_cellmath__24_0_I999 (.Y(N2429), .A(N2511));
OAI22XL inst_cellmath__24_0_I1000 (.Y(N3641), .A0(N2429), .A1(N2320), .B0(N3305), .B1(N2963));
INVXL inst_cellmath__24_0_I1001 (.Y(N3110), .A(N2853));
OAI22XL inst_cellmath__24_0_I1002 (.Y(N2774), .A0(N3110), .A1(N2320), .B0(N2429), .B1(N2963));
INVXL inst_cellmath__24_0_I1003 (.Y(N2230), .A(N3186));
OAI22XL inst_cellmath__24_0_I1004 (.Y(N3448), .A0(N2230), .A1(N2320), .B0(N3110), .B1(N2963));
INVXL inst_cellmath__24_0_I1005 (.Y(N2914), .A(N3513));
OAI22XL inst_cellmath__24_0_I1006 (.Y(N2576), .A0(N2914), .A1(N2320), .B0(N2230), .B1(N2963));
INVXL inst_cellmath__24_0_I1007 (.Y(N3581), .A(N2308));
OAI22XL inst_cellmath__24_0_I1008 (.Y(N3245), .A0(N3581), .A1(N2320), .B0(N2914), .B1(N2963));
INVXL inst_cellmath__24_0_I1009 (.Y(N2714), .A(N2653));
OAI22XL inst_cellmath__24_0_I1010 (.Y(N2372), .A0(N2714), .A1(N2320), .B0(N3581), .B1(N2963));
INVXL inst_cellmath__24_0_I1011 (.Y(N3395), .A(N2987));
OAI22XL inst_cellmath__24_0_I1012 (.Y(N3050), .A0(N3395), .A1(N2320), .B0(N2714), .B1(N2963));
INVXL inst_cellmath__24_0_I1013 (.Y(N2516), .A(N3329));
OAI22XL inst_cellmath__24_0_I1014 (.Y(N2175), .A0(N2516), .A1(N2320), .B0(N3395), .B1(N2963));
INVXL inst_cellmath__24_0_I1015 (.Y(N3190), .A(N3660));
OAI22XL inst_cellmath__24_0_I1016 (.Y(N2857), .A0(N3190), .A1(N2320), .B0(N2516), .B1(N2963));
INVXL inst_cellmath__24_0_I1017 (.Y(N2313), .A(N2452));
OAI22XL inst_cellmath__24_0_I1018 (.Y(N3518), .A0(N2313), .A1(N2320), .B0(N3190), .B1(N2963));
INVXL inst_cellmath__24_0_I1019 (.Y(N2990), .A(N2799));
OAI22XL inst_cellmath__24_0_I1020 (.Y(N2657), .A0(N2990), .A1(N2320), .B0(N2313), .B1(N2963));
INVXL inst_cellmath__24_0_I1021 (.Y(N3664), .A(N3134));
OAI22XL inst_cellmath__24_0_I1022 (.Y(N3333), .A0(N3664), .A1(N2320), .B0(N2990), .B1(N2963));
NOR2XL inst_cellmath__24_0_I1023 (.Y(N2454), .A(N3664), .B(N2963));
INVXL inst_cellmath__24_0_I1024 (.Y(N3136), .A(N2320));
NAND2XL inst_cellmath__24_0_I1025 (.Y(N2938), .A(N2320), .B(N2963));
AO21XL inst_cellmath__24_0_I1026 (.Y(N2677), .A0(N2357), .A1(N2935), .B0(N3272));
AO21XL inst_cellmath__24_0_I1027 (.Y(N3012), .A0(N8302), .A1(N2620), .B0(N2959));
AO21XL inst_cellmath__24_0_I1028 (.Y(N3350), .A0(N8310), .A1(N2302), .B0(N2645));
AO21XL inst_cellmath__24_0_I1029 (.Y(N3680), .A0(N8327), .A1(N3175), .B0(N2332));
AO21XL inst_cellmath__24_0_I1030 (.Y(N2473), .A0(N8335), .A1(N3114), .B0(N3564));
AO21XL inst_cellmath__24_0_I1031 (.Y(N2817), .A0(N8342), .A1(N3048), .B0(N3258));
AO21XL inst_cellmath__24_0_I1032 (.Y(N3152), .A0(N2646), .A1(N2981), .B0(N2947));
AO21XL inst_cellmath__24_0_I1033 (.Y(N3481), .A0(N8358), .A1(N2923), .B0(N2352));
AO21XL inst_cellmath__24_0_I1034 (.Y(N2273), .A0(N2519), .A1(N2860), .B0(N3583));
AO21XL inst_cellmath__24_0_I1035 (.Y(N2615), .A0(N2450), .A1(N2659), .B0(N2993));
AO21XL inst_cellmath__24_0_I1036 (.Y(N2955), .A0(N2385), .A1(N3609), .B0(N2395));
ADDHX1 inst_cellmath__24_0_I1037 (.CO(N3626), .S(N3290), .A(N3446), .B(N3647));
ADDHX1 inst_cellmath__24_0_I1038 (.CO(N2759), .S(N2412), .A(N2781), .B(N2913));
ADDHX1 inst_cellmath__24_0_I1039 (.CO(N3436), .S(N3095), .A(N3385), .B(N3452));
ADDFX1 inst_cellmath__24_0_I1040 (.CO(N2561), .S(N2215), .A(N2166), .B(N3582), .CI(N2759));
ADDHX1 inst_cellmath__24_0_I1041 (.CO(N3231), .S(N2899), .A(N2584), .B(N2715));
ADDFX1 inst_cellmath__24_0_I1042 (.CO(N2362), .S(N3569), .A(N3436), .B(N2850), .CI(N2899));
ADDHX1 inst_cellmath__24_0_I1043 (.CO(N3037), .S(N2700), .A(N3317), .B(N3253));
ADDFX1 inst_cellmath__24_0_I1044 (.CO(N2499), .S(N3260), .A(N3510), .B(N3396), .CI(N3650));
ADDFX1 inst_cellmath__24_0_I1045 (.CO(N2161), .S(N3377), .A(N3231), .B(N2700), .CI(N3260));
ADDHX1 inst_cellmath__24_0_I1046 (.CO(N3174), .S(N2846), .A(N2378), .B(N2517));
ADDFX1 inst_cellmath__24_0_I1047 (.CO(N3319), .S(N2977), .A(N2786), .B(N2649), .CI(N3037));
ADDFX1 inst_cellmath__24_0_I1048 (.CO(N2439), .S(N3649), .A(N2499), .B(N2846), .CI(N2977));
ADDHX1 inst_cellmath__24_0_I1049 (.CO(N3121), .S(N2788), .A(N3251), .B(N3054));
ADDFX1 inst_cellmath__24_0_I1050 (.CO(N2245), .S(N3456), .A(N3324), .B(N3188), .CI(N3457));
ADDFX1 inst_cellmath__24_0_I1051 (.CO(N3263), .S(N3001), .A(N3174), .B(N3586), .CI(N2788));
ADDFX1 inst_cellmath__24_0_I1052 (.CO(N2926), .S(N2588), .A(N3319), .B(N3456), .CI(N3001));
ADDHX1 inst_cellmath__24_0_I1053 (.CO(N2382), .S(N3592), .A(N2180), .B(N2314));
ADDFX1 inst_cellmath__24_0_I1054 (.CO(N3061), .S(N2727), .A(N2589), .B(N2448), .CI(N2718));
ADDFX1 inst_cellmath__24_0_I1055 (.CO(N3202), .S(N2868), .A(N3592), .B(N3121), .CI(N2245));
ADDFX1 inst_cellmath__24_0_I1056 (.CO(N2327), .S(N3531), .A(N2727), .B(N3263), .CI(N2868));
ADDHX1 inst_cellmath__24_0_I1057 (.CO(N3002), .S(N2671), .A(N3185), .B(N2863));
ADDFX1 inst_cellmath__24_0_I1058 (.CO(N2466), .S(N2752), .A(N3129), .B(N2991), .CI(N3261));
ADDFX1 inst_cellmath__24_0_I1059 (.CO(N3674), .S(N3344), .A(N3061), .B(N2671), .CI(N2752));
ADDFX1 inst_cellmath__24_0_I1060 (.CO(N2608), .S(N2265), .A(N3515), .B(N3400), .CI(N2382));
ADDFX1 inst_cellmath__24_0_I1061 (.CO(N3283), .S(N2948), .A(N3202), .B(N2265), .CI(N3344));
ADDHX1 inst_cellmath__24_0_I1062 (.CO(N2407), .S(N3619), .A(N3525), .B(N3662));
ADDFX1 inst_cellmath__24_0_I1063 (.CO(N3429), .S(N2491), .A(N2383), .B(N2249), .CI(N2520));
ADDFX1 inst_cellmath__24_0_I1064 (.CO(N3088), .S(N2753), .A(N3619), .B(N2466), .CI(N2491));
ADDFX1 inst_cellmath__24_0_I1065 (.CO(N3557), .S(N3225), .A(N3002), .B(N2652), .CI(N2608));
ADDFX1 inst_cellmath__24_0_I1066 (.CO(N2694), .S(N2355), .A(N3225), .B(N3674), .CI(N2753));
ADDHX1 inst_cellmath__24_0_I1067 (.CO(N3369), .S(N3029), .A(N3126), .B(N2664));
ADDFX1 inst_cellmath__24_0_I1068 (.CO(N2492), .S(N2155), .A(N2932), .B(N2802), .CI(N3062));
ADDFX1 inst_cellmath__24_0_I1069 (.CO(N3499), .S(N2235), .A(N3331), .B(N3193), .CI(N3460));
ADDFX1 inst_cellmath__24_0_I1070 (.CO(N3169), .S(N2839), .A(N3029), .B(N3429), .CI(N2235));
ADDFX1 inst_cellmath__24_0_I1071 (.CO(N3644), .S(N3311), .A(N2155), .B(N2407), .CI(N3557));
ADDFX1 inst_cellmath__24_0_I1072 (.CO(N2780), .S(N2433), .A(N2839), .B(N3088), .CI(N3311));
ADDHX1 inst_cellmath__24_0_I1073 (.CO(N3450), .S(N3113), .A(N3341), .B(N3466));
ADDFX1 inst_cellmath__24_0_I1074 (.CO(N2581), .S(N2236), .A(N2185), .B(N3600), .CI(N2318));
ADDFX1 inst_cellmath__24_0_I1075 (.CO(N2719), .S(N2374), .A(N2592), .B(N2453), .CI(N3369));
ADDFX1 inst_cellmath__24_0_I1076 (.CO(N3399), .S(N3052), .A(N3499), .B(N3113), .CI(N2492));
ADDFX1 inst_cellmath__24_0_I1077 (.CO(N3523), .S(N3194), .A(N2374), .B(N2236), .CI(N3169));
ADDFX1 inst_cellmath__24_0_I1078 (.CO(N2663), .S(N2317), .A(N3644), .B(N3052), .CI(N3194));
ADDHX1 inst_cellmath__24_0_I1079 (.CO(N3338), .S(N2995), .A(N3058), .B(N2461));
ADDFX1 inst_cellmath__24_0_I1080 (.CO(N2805), .S(N3522), .A(N2733), .B(N2598), .CI(N2869));
ADDFX1 inst_cellmath__24_0_I1081 (.CO(N2459), .S(N3668), .A(N2581), .B(N2995), .CI(N3522));
ADDFX1 inst_cellmath__24_0_I1082 (.CO(N2260), .S(N3277), .A(N3133), .B(N2996), .CI(N3267));
ADDFX1 inst_cellmath__24_0_I1083 (.CO(N3469), .S(N3142), .A(N3403), .B(N3450), .CI(N3277));
ADDFX1 inst_cellmath__24_0_I1084 (.CO(N2398), .S(N3614), .A(N3399), .B(N2719), .CI(N3668));
ADDFX1 inst_cellmath__24_0_I1085 (.CO(N3082), .S(N2744), .A(N3523), .B(N3142), .CI(N3614));
ADDHX1 inst_cellmath__24_0_I1086 (.CO(N2200), .S(N3421), .A(N3143), .B(N3275));
ADDFX1 inst_cellmath__24_0_I1087 (.CO(N3218), .S(N3022), .A(N3532), .B(N3411), .CI(N3667));
ADDFX1 inst_cellmath__24_0_I1088 (.CO(N2885), .S(N2547), .A(N2260), .B(N2805), .CI(N3022));
ADDFX1 inst_cellmath__24_0_I1089 (.CO(N2687), .S(N2771), .A(N2387), .B(N2255), .CI(N2523));
ADDFX1 inst_cellmath__24_0_I1090 (.CO(N2347), .S(N3552), .A(N3338), .B(N3421), .CI(N2771));
ADDFX1 inst_cellmath__24_0_I1091 (.CO(N2832), .S(N2485), .A(N3469), .B(N2459), .CI(N2547));
ADDFX1 inst_cellmath__24_0_I1092 (.CO(N3494), .S(N3165), .A(N2398), .B(N3552), .CI(N2485));
ADDHX1 inst_cellmath__24_0_I1093 (.CO(N2628), .S(N2286), .A(N2994), .B(N2263));
ADDFX1 inst_cellmath__24_0_I1094 (.CO(N3304), .S(N2966), .A(N2535), .B(N2394), .CI(N2669));
ADDFX1 inst_cellmath__24_0_I1095 (.CO(N2773), .S(N2512), .A(N2937), .B(N2806), .CI(N3065));
ADDFX1 inst_cellmath__24_0_I1096 (.CO(N2427), .S(N3638), .A(N2687), .B(N3218), .CI(N2512));
ADDFX1 inst_cellmath__24_0_I1097 (.CO(N2912), .S(N2575), .A(N3200), .B(N3336), .CI(N2200));
ADDFX1 inst_cellmath__24_0_I1098 (.CO(N3579), .S(N3244), .A(N2966), .B(N2286), .CI(N2575));
ADDFX1 inst_cellmath__24_0_I1099 (.CO(N2172), .S(N3392), .A(N2347), .B(N2885), .CI(N3244));
ADDFX1 inst_cellmath__24_0_I1100 (.CO(N2854), .S(N2513), .A(N2832), .B(N3638), .CI(N3392));
ADDHX1 inst_cellmath__24_0_I1101 (.CO(N3514), .S(N3187), .A(N2943), .B(N3074));
ADDFX1 inst_cellmath__24_0_I1102 (.CO(N2654), .S(N2310), .A(N3345), .B(N3207), .CI(N3470));
ADDFX1 inst_cellmath__24_0_I1103 (.CO(N3661), .S(N2253), .A(N2189), .B(N3607), .CI(N2323));
ADDFX1 inst_cellmath__24_0_I1104 (.CO(N3330), .S(N2988), .A(N3304), .B(N2773), .CI(N2253));
ADDFX1 inst_cellmath__24_0_I1105 (.CO(N2254), .S(N3464), .A(N2628), .B(N2458), .CI(N3187));
ADDFX1 inst_cellmath__24_0_I1106 (.CO(N2936), .S(N2597), .A(N2310), .B(N2912), .CI(N3464));
ADDFX1 inst_cellmath__24_0_I1107 (.CO(N3073), .S(N2737), .A(N3579), .B(N2427), .CI(N2988));
ADDFX1 inst_cellmath__24_0_I1108 (.CO(N2193), .S(N3415), .A(N2172), .B(N2597), .CI(N2737));
ADDHX1 inst_cellmath__24_0_I1109 (.CO(N2878), .S(N2540), .A(N2933), .B(N3615));
ADDFX1 inst_cellmath__24_0_I1110 (.CO(N2340), .S(N3541), .A(N2196), .B(N2467), .CI(N2335));
ADDFX1 inst_cellmath__24_0_I1111 (.CO(N3544), .S(N3212), .A(N2654), .B(N3661), .CI(N3541));
ADDFX1 inst_cellmath__24_0_I1112 (.CO(N3357), .S(N3295), .A(N2738), .B(N2603), .CI(N2873));
ADDFX1 inst_cellmath__24_0_I1113 (.CO(N3018), .S(N2682), .A(N3514), .B(N2540), .CI(N3295));
ADDFX1 inst_cellmath__24_0_I1114 (.CO(N3487), .S(N3159), .A(N3137), .B(N2999), .CI(N3271));
ADDFX1 inst_cellmath__24_0_I1115 (.CO(N2622), .S(N2278), .A(N2254), .B(N3159), .CI(N3330));
ADDFX1 inst_cellmath__24_0_I1116 (.CO(N3632), .S(N3040), .A(N3212), .B(N2936), .CI(N2682));
ADDFX1 inst_cellmath__24_0_I1117 (.CO(N3296), .S(N2960), .A(N3073), .B(N2278), .CI(N3040));
ADDHX1 inst_cellmath__24_0_I1118 (.CO(N2764), .S(N2420), .A(N2749), .B(N2880));
ADDFX1 inst_cellmath__24_0_I1119 (.CO(N2221), .S(N2791), .A(N3147), .B(N3010), .CI(N3278));
ADDFX1 inst_cellmath__24_0_I1120 (.CO(N3441), .S(N3102), .A(N3487), .B(N2340), .CI(N2791));
ADDFX1 inst_cellmath__24_0_I1121 (.CO(N3236), .S(N2532), .A(N3535), .B(N3416), .CI(N3672));
ADDFX1 inst_cellmath__24_0_I1122 (.CO(N2905), .S(N2566), .A(N2420), .B(N3357), .CI(N2532));
ADDFX1 inst_cellmath__24_0_I1123 (.CO(N3384), .S(N3042), .A(N2392), .B(N2259), .CI(N2878));
ADDFX1 inst_cellmath__24_0_I1124 (.CO(N2504), .S(N2164), .A(N3544), .B(N3042), .CI(N3018));
ADDFX1 inst_cellmath__24_0_I1125 (.CO(N3508), .S(N2271), .A(N2566), .B(N3102), .CI(N2622));
ADDFX1 inst_cellmath__24_0_I1126 (.CO(N3182), .S(N2849), .A(N2164), .B(N3632), .CI(N2271));
ADDHX1 inst_cellmath__24_0_I1127 (.CO(N2648), .S(N2303), .A(N2871), .B(N3424));
ADDFX1 inst_cellmath__24_0_I1128 (.CO(N3323), .S(N2980), .A(N3681), .B(N3545), .CI(N2266));
ADDFX1 inst_cellmath__24_0_I1129 (.CO(N2794), .S(N3563), .A(N2539), .B(N2399), .CI(N2675));
ADDFX1 inst_cellmath__24_0_I1130 (.CO(N2443), .S(N3654), .A(N3236), .B(N2221), .CI(N3563));
ADDFX1 inst_cellmath__24_0_I1131 (.CO(N2247), .S(N3315), .A(N2941), .B(N2811), .CI(N3070));
ADDFX1 inst_cellmath__24_0_I1132 (.CO(N3459), .S(N3128), .A(N2764), .B(N2303), .CI(N3315));
ADDFX1 inst_cellmath__24_0_I1133 (.CO(N2386), .S(N3599), .A(N3384), .B(N3204), .CI(N2980));
ADDFX1 inst_cellmath__24_0_I1134 (.CO(N3066), .S(N2730), .A(N2905), .B(N3441), .CI(N3599));
ADDFX1 inst_cellmath__24_0_I1135 (.CO(N2534), .S(N3056), .A(N3128), .B(N3654), .CI(N2504));
ADDFX1 inst_cellmath__24_0_I1136 (.CO(N2188), .S(N3409), .A(N2730), .B(N3508), .CI(N3056));
ADDHX1 inst_cellmath__24_0_I1137 (.CO(N3205), .S(N2872), .A(N2548), .B(N2684));
ADDFX1 inst_cellmath__24_0_I1138 (.CO(N2333), .S(N3536), .A(N2949), .B(N2818), .CI(N3080));
ADDFX1 inst_cellmath__24_0_I1139 (.CO(N3347), .S(N2809), .A(N3348), .B(N3213), .CI(N3472));
ADDFX1 inst_cellmath__24_0_I1140 (.CO(N3009), .S(N2674), .A(N3323), .B(N2794), .CI(N2809));
ADDFX1 inst_cellmath__24_0_I1141 (.CO(N2815), .S(N2551), .A(N2192), .B(N3612), .CI(N2330));
ADDFX1 inst_cellmath__24_0_I1142 (.CO(N2471), .S(N3677), .A(N2872), .B(N2247), .CI(N2551));
ADDFX1 inst_cellmath__24_0_I1143 (.CO(N2953), .S(N2612), .A(N3536), .B(N2648), .CI(N2386));
ADDFX1 inst_cellmath__24_0_I1144 (.CO(N3624), .S(N3288), .A(N3459), .B(N2443), .CI(N3677));
ADDFX1 inst_cellmath__24_0_I1145 (.CO(N2213), .S(N3433), .A(N3066), .B(N2674), .CI(N2612));
ADDFX1 inst_cellmath__24_0_I1146 (.CO(N2896), .S(N2558), .A(N2534), .B(N3288), .CI(N3433));
ADDHX1 inst_cellmath__24_0_I1147 (.CO(N3566), .S(N3228), .A(N2807), .B(N2400));
ADDFX1 inst_cellmath__24_0_I1148 (.CO(N3034), .S(N2290), .A(N3361), .B(N3221), .CI(N3480));
ADDFX1 inst_cellmath__24_0_I1149 (.CO(N2698), .S(N2360), .A(N2333), .B(N3347), .CI(N2290));
ADDFX1 inst_cellmath__24_0_I1150 (.CO(N2496), .S(N3584), .A(N2201), .B(N3620), .CI(N2341));
ADDFX1 inst_cellmath__24_0_I1151 (.CO(N2158), .S(N3375), .A(N3205), .B(N2815), .CI(N3584));
ADDFX1 inst_cellmath__24_0_I1152 (.CO(N2638), .S(N2297), .A(N2470), .B(N3005), .CI(N2606));
ADDFX1 inst_cellmath__24_0_I1153 (.CO(N3316), .S(N2975), .A(N2877), .B(N2743), .CI(N3228));
ADDFX1 inst_cellmath__24_0_I1154 (.CO(N3454), .S(N3119), .A(N2975), .B(N2297), .CI(N2471));
ADDFX1 inst_cellmath__24_0_I1155 (.CO(N2585), .S(N2241), .A(N3375), .B(N3009), .CI(N2360));
ADDFX1 inst_cellmath__24_0_I1156 (.CO(N3590), .S(N3335), .A(N3119), .B(N2953), .CI(N3624));
ADDFX1 inst_cellmath__24_0_I1157 (.CO(N3259), .S(N2922), .A(N2241), .B(N2213), .CI(N3335));
ADDHX1 inst_cellmath__24_0_I1158 (.CO(N2724), .S(N2379), .A(N3085), .B(N2350));
ADDFX1 inst_cellmath__24_0_I1159 (.CO(N2183), .S(N3076), .A(N3566), .B(N2479), .CI(N2616));
ADDFX1 inst_cellmath__24_0_I1160 (.CO(N3402), .S(N3057), .A(N2638), .B(N3034), .CI(N3076));
ADDFX1 inst_cellmath__24_0_I1161 (.CO(N3199), .S(N2828), .A(N2886), .B(N2754), .CI(N3016));
ADDFX1 inst_cellmath__24_0_I1162 (.CO(N2864), .S(N2525), .A(N3316), .B(N2496), .CI(N2828));
ADDFX1 inst_cellmath__24_0_I1163 (.CO(N2666), .S(N2570), .A(N3282), .B(N3151), .CI(N3419));
ADDFX1 inst_cellmath__24_0_I1164 (.CO(N2322), .S(N3530), .A(N3538), .B(N2379), .CI(N2570));
ADDFX1 inst_cellmath__24_0_I1165 (.CO(N2810), .S(N2465), .A(N2698), .B(N3676), .CI(N2158));
ADDFX1 inst_cellmath__24_0_I1166 (.CO(N3473), .S(N3145), .A(N3530), .B(N3057), .CI(N2525));
ADDFX1 inst_cellmath__24_0_I1167 (.CO(N3617), .S(N3281), .A(N2465), .B(N3454), .CI(N2585));
ADDFX1 inst_cellmath__24_0_I1168 (.CO(N2750), .S(N2404), .A(N3590), .B(N3145), .CI(N3281));
ADDFX1 inst_cellmath__24_0_I1169 (.CO(N3427), .S(N3086), .A(N2203), .B(N2748), .CI(N3162));
ADDFX1 inst_cellmath__24_0_I1170 (.CO(N2891), .S(N2306), .A(N3024), .B(N3291), .CI(N3428));
ADDFX1 inst_cellmath__24_0_I1171 (.CO(N2553), .S(N2205), .A(N2666), .B(N3199), .CI(N2306));
ADDFX1 inst_cellmath__24_0_I1172 (.CO(N2353), .S(N3602), .A(N3686), .B(N3551), .CI(N2272));
ADDFX1 inst_cellmath__24_0_I1173 (.CO(N3555), .S(N3222), .A(N2724), .B(N2183), .CI(N3602));
ADDFX1 inst_cellmath__24_0_I1174 (.CO(N3367), .S(N3353), .A(N2545), .B(N2403), .CI(N2680));
ADDFX1 inst_cellmath__24_0_I1175 (.CO(N3027), .S(N2692), .A(N3086), .B(N2814), .CI(N3353));
ADDFX1 inst_cellmath__24_0_I1176 (.CO(N2837), .S(N3097), .A(N2864), .B(N3402), .CI(N2322));
ADDFX1 inst_cellmath__24_0_I1177 (.CO(N2489), .S(N2152), .A(N3222), .B(N2810), .CI(N3097));
ADDFX1 inst_cellmath__24_0_I1178 (.CO(N2971), .S(N2633), .A(N2692), .B(N2205), .CI(N3473));
ADDFX1 inst_cellmath__24_0_I1179 (.CO(N3642), .S(N3309), .A(N2633), .B(N3617), .CI(N2152));
INVXL inst_cellmath__24_0_I1180 (.Y(N2641), .A(N3423));
ADDFX1 inst_cellmath__24_0_I1181 (.CO(N2778), .S(N2431), .A(N2282), .B(N2887), .CI(N2641));
ADDFX1 inst_cellmath__24_0_I1182 (.CO(N2915), .S(N2789), .A(N2555), .B(N2411), .CI(N2688));
ADDFX1 inst_cellmath__24_0_I1183 (.CO(N2579), .S(N2234), .A(N3367), .B(N2353), .CI(N2789));
ADDFX1 inst_cellmath__24_0_I1184 (.CO(N2373), .S(N2528), .A(N2952), .B(N2822), .CI(N3087));
ADDFX1 inst_cellmath__24_0_I1185 (.CO(N3585), .S(N3249), .A(N3427), .B(N2891), .CI(N2528));
ADDFX1 inst_cellmath__24_0_I1186 (.CO(N2518), .S(N2178), .A(N3355), .B(N3217), .CI(N3476));
ADDFX1 inst_cellmath__24_0_I1187 (.CO(N3192), .S(N2859), .A(N2178), .B(N2677), .CI(N2431));
ADDFX1 inst_cellmath__24_0_I1188 (.CO(N2661), .S(N2268), .A(N3555), .B(N2553), .CI(N3027));
ADDFX1 inst_cellmath__24_0_I1189 (.CO(N2316), .S(N3521), .A(N2234), .B(N2837), .CI(N2268));
ADDFX1 inst_cellmath__24_0_I1190 (.CO(N2803), .S(N2457), .A(N3249), .B(N2859), .CI(N2489));
ADDFX1 inst_cellmath__24_0_I1191 (.CO(N3467), .S(N3139), .A(N3521), .B(N2971), .CI(N2457));
INVXL inst_cellmath__24_0_I1192 (.Y(N3370), .A(N2550));
ADDFX1 inst_cellmath__24_0_I1193 (.CO(N2602), .S(N2258), .A(N3554), .B(N3423), .CI(N3370));
ADDFX1 inst_cellmath__24_0_I1194 (.CO(N2742), .S(N3500), .A(N2962), .B(N3096), .CI(N3226));
ADDFX1 inst_cellmath__24_0_I1195 (.CO(N2396), .S(N3611), .A(N2518), .B(N2778), .CI(N3500));
ADDFX1 inst_cellmath__24_0_I1196 (.CO(N2198), .S(N3252), .A(N3485), .B(N3363), .CI(N3625));
ADDFX1 inst_cellmath__24_0_I1197 (.CO(N3420), .S(N3078), .A(N2373), .B(N2915), .CI(N3252));
ADDFX1 inst_cellmath__24_0_I1198 (.CO(N3216), .S(N2997), .A(N2345), .B(N2206), .CI(N2474));
ADDFX1 inst_cellmath__24_0_I1199 (.CO(N2883), .S(N2544), .A(N2611), .B(N2258), .CI(N2997));
ADDFX1 inst_cellmath__24_0_I1200 (.CO(N2685), .S(N2746), .A(N3192), .B(N2579), .CI(N3585));
ADDFX1 inst_cellmath__24_0_I1201 (.CO(N2346), .S(N3549), .A(N3078), .B(N2661), .CI(N2746));
ADDFX1 inst_cellmath__24_0_I1202 (.CO(N2831), .S(N2482), .A(N2544), .B(N3611), .CI(N2316));
ADDFX1 inst_cellmath__24_0_I1203 (.CO(N3491), .S(N3163), .A(N2803), .B(N3549), .CI(N2482));
ADDFX1 inst_cellmath__24_0_I1204 (.CO(N2625), .S(N2285), .A(N2550), .B(N3220), .CI(N2690));
ADDFX1 inst_cellmath__24_0_I1205 (.CO(N3636), .S(N2486), .A(N2354), .B(N2216), .CI(N2484));
ADDFX1 inst_cellmath__24_0_I1206 (.CO(N3302), .S(N2964), .A(N3216), .B(N2198), .CI(N2486));
ADDFX1 inst_cellmath__24_0_I1207 (.CO(N3106), .S(N2229), .A(N2758), .B(N2623), .CI(N2890));
ADDFX1 inst_cellmath__24_0_I1208 (.CO(N2770), .S(N2424), .A(N2602), .B(N2742), .CI(N2229));
ADDFX1 inst_cellmath__24_0_I1209 (.CO(N2571), .S(N3517), .A(N3156), .B(N3021), .CI(N3287));
ADDFX1 inst_cellmath__24_0_I1210 (.CO(N2227), .S(N3443), .A(N3012), .B(N2285), .CI(N3517));
ADDFX1 inst_cellmath__24_0_I1211 (.CO(N3575), .S(N3274), .A(N3420), .B(N2396), .CI(N2883));
ADDFX1 inst_cellmath__24_0_I1212 (.CO(N3242), .S(N2909), .A(N2964), .B(N2685), .CI(N3274));
ADDFX1 inst_cellmath__24_0_I1213 (.CO(N2170), .S(N3389), .A(N3443), .B(N2424), .CI(N2346));
ADDFX1 inst_cellmath__24_0_I1214 (.CO(N2852), .S(N2508), .A(N2831), .B(N2909), .CI(N3389));
INVXL inst_cellmath__24_0_I1215 (.Y(N2824), .A(N2349));
ADDFX1 inst_cellmath__24_0_I1216 (.CO(N3511), .S(N3184), .A(N3030), .B(N3364), .CI(N2824));
ADDFX1 inst_cellmath__24_0_I1217 (.CO(N3328), .S(N2986), .A(N3297), .B(N3166), .CI(N2897));
ADDFX1 inst_cellmath__24_0_I1218 (.CO(N2798), .S(N2961), .A(N3556), .B(N3432), .CI(N3689));
ADDFX1 inst_cellmath__24_0_I1219 (.CO(N2449), .S(N3658), .A(N3106), .B(N3636), .CI(N2961));
ADDFX1 inst_cellmath__24_0_I1220 (.CO(N2252), .S(N2708), .A(N2408), .B(N2277), .CI(N2625));
ADDFX1 inst_cellmath__24_0_I1221 (.CO(N3463), .S(N3132), .A(N2986), .B(N3184), .CI(N2708));
ADDFX1 inst_cellmath__24_0_I1222 (.CO(N2391), .S(N3605), .A(N2227), .B(N2571), .CI(N3302));
ADDFX1 inst_cellmath__24_0_I1223 (.CO(N3071), .S(N2735), .A(N3658), .B(N2770), .CI(N3132));
ADDFX1 inst_cellmath__24_0_I1224 (.CO(N3210), .S(N2876), .A(N3605), .B(N3575), .CI(N2735));
ADDFX1 inst_cellmath__24_0_I1225 (.CO(N2337), .S(N3540), .A(N2170), .B(N3242), .CI(N2876));
ADDFX1 inst_cellmath__24_0_I1226 (.CO(N3354), .S(N2446), .A(N2349), .B(N3026), .CI(N2487));
ADDFX1 inst_cellmath__24_0_I1227 (.CO(N3015), .S(N2679), .A(N2156), .B(N3350), .CI(N2446));
ADDFX1 inst_cellmath__24_0_I1228 (.CO(N2819), .S(N2190), .A(N2418), .B(N2287), .CI(N2559));
ADDFX1 inst_cellmath__24_0_I1229 (.CO(N2475), .S(N3683), .A(N3328), .B(N3511), .CI(N2190));
ADDFX1 inst_cellmath__24_0_I1230 (.CO(N2276), .S(N3479), .A(N2829), .B(N2693), .CI(N2956));
ADDFX1 inst_cellmath__24_0_I1231 (.CO(N3484), .S(N3155), .A(N3093), .B(N2798), .CI(N3479));
ADDFX1 inst_cellmath__24_0_I1232 (.CO(N2416), .S(N3629), .A(N2679), .B(N2252), .CI(N2449));
ADDFX1 inst_cellmath__24_0_I1233 (.CO(N3098), .S(N2763), .A(N3155), .B(N3463), .CI(N3683));
ADDFX1 inst_cellmath__24_0_I1234 (.CO(N2563), .S(N3230), .A(N3629), .B(N2391), .CI(N3071));
ADDFX1 inst_cellmath__24_0_I1235 (.CO(N2220), .S(N3437), .A(N2763), .B(N3210), .CI(N3230));
INVXL inst_cellmath__24_0_I1236 (.Y(N2785), .A(N2150));
ADDFX1 inst_cellmath__24_0_I1237 (.CO(N3235), .S(N2901), .A(N2967), .B(N3167), .CI(N2785));
ADDFX1 inst_cellmath__24_0_I1238 (.CO(N3380), .S(N2924), .A(N2838), .B(N3103), .CI(N3229));
ADDFX1 inst_cellmath__24_0_I1239 (.CO(N3038), .S(N2705), .A(N2276), .B(N2819), .CI(N2924));
ADDFX1 inst_cellmath__24_0_I1240 (.CO(N3506), .S(N3179), .A(N3492), .B(N3366), .CI(N3630));
ADDFX1 inst_cellmath__24_0_I1241 (.CO(N2644), .S(N2299), .A(N3354), .B(N2210), .CI(N3179));
ADDFX1 inst_cellmath__24_0_I1242 (.CO(N2790), .S(N2441), .A(N3015), .B(N2901), .CI(N3484));
ADDFX1 inst_cellmath__24_0_I1243 (.CO(N3458), .S(N3125), .A(N2299), .B(N2475), .CI(N2705));
ADDFX1 inst_cellmath__24_0_I1244 (.CO(N3596), .S(N3265), .A(N2441), .B(N2416), .CI(N3098));
ADDFX1 inst_cellmath__24_0_I1245 (.CO(N2729), .S(N2384), .A(N2563), .B(N3125), .CI(N3265));
ADDFX1 inst_cellmath__24_0_I1246 (.CO(N3408), .S(N3064), .A(N2150), .B(N2835), .CI(N2288));
ADDFX1 inst_cellmath__24_0_I1247 (.CO(N2870), .S(N2668), .A(N2222), .B(N3639), .CI(N2359));
ADDFX1 inst_cellmath__24_0_I1248 (.CO(N2530), .S(N2187), .A(N3506), .B(N3235), .CI(N2668));
ADDFX1 inst_cellmath__24_0_I1249 (.CO(N2329), .S(N2405), .A(N2626), .B(N2490), .CI(N2762));
ADDFX1 inst_cellmath__24_0_I1250 (.CO(N3534), .S(N3203), .A(N3064), .B(N3380), .CI(N2405));
ADDFX1 inst_cellmath__24_0_I1251 (.CO(N2469), .S(N3675), .A(N3680), .B(N2893), .CI(N3038));
ADDFX1 inst_cellmath__24_0_I1252 (.CO(N3149), .S(N2813), .A(N3203), .B(N2644), .CI(N2187));
ADDFX1 inst_cellmath__24_0_I1253 (.CO(N2610), .S(N2154), .A(N3675), .B(N2790), .CI(N3458));
ADDFX1 inst_cellmath__24_0_I1254 (.CO(N2269), .S(N3477), .A(N2813), .B(N3596), .CI(N2154));
INVXL inst_cellmath__24_0_I1255 (.Y(N3250), .A(N3497));
ADDFX1 inst_cellmath__24_0_I1256 (.CO(N3286), .S(N2951), .A(N2903), .B(N2970), .CI(N3250));
ADDFX1 inst_cellmath__24_0_I1257 (.CO(N3092), .S(N2756), .A(N3168), .B(N3035), .CI(N2772));
ADDFX1 inst_cellmath__24_0_I1258 (.CO(N2556), .S(N3398), .A(N3438), .B(N3300), .CI(N3562));
ADDFX1 inst_cellmath__24_0_I1259 (.CO(N2209), .S(N3431), .A(N2329), .B(N2870), .CI(N3398));
ADDFX1 inst_cellmath__24_0_I1260 (.CO(N2696), .S(N2358), .A(N2756), .B(N3408), .CI(N2951));
ADDFX1 inst_cellmath__24_0_I1261 (.CO(N3372), .S(N3031), .A(N3534), .B(N2530), .CI(N2358));
ADDFX1 inst_cellmath__24_0_I1262 (.CO(N3501), .S(N3171), .A(N2469), .B(N3431), .CI(N3149));
ADDFX1 inst_cellmath__24_0_I1263 (.CO(N2637), .S(N2293), .A(N2610), .B(N3031), .CI(N3171));
ADDFX1 inst_cellmath__24_0_I1264 (.CO(N3648), .S(N3140), .A(N3497), .B(N2631), .CI(N3641));
ADDFX1 inst_cellmath__24_0_I1265 (.CO(N3313), .S(N2973), .A(N3573), .B(N2473), .CI(N3140));
ADDFX1 inst_cellmath__24_0_I1266 (.CO(N3117), .S(N2884), .A(N2291), .B(N2159), .CI(N2425));
ADDFX1 inst_cellmath__24_0_I1267 (.CO(N2782), .S(N2435), .A(N3092), .B(N3286), .CI(N2884));
ADDFX1 inst_cellmath__24_0_I1268 (.CO(N3255), .S(N2918), .A(N2697), .B(N2564), .CI(N2556));
ADDFX1 inst_cellmath__24_0_I1269 (.CO(N2376), .S(N3589), .A(N2918), .B(N2973), .CI(N2209));
ADDFX1 inst_cellmath__24_0_I1270 (.CO(N2522), .S(N2181), .A(N2435), .B(N2696), .CI(N3589));
ADDFX1 inst_cellmath__24_0_I1271 (.CO(N3196), .S(N2862), .A(N3501), .B(N3372), .CI(N2181));
INVXL inst_cellmath__24_0_I1272 (.Y(N2426), .A(N3305));
ADDFX1 inst_cellmath__24_0_I1273 (.CO(N2319), .S(N3527), .A(N2843), .B(N2774), .CI(N2426));
ADDFX1 inst_cellmath__24_0_I1274 (.CO(N2462), .S(N2574), .A(N2706), .B(N2972), .CI(N3107));
ADDFX1 inst_cellmath__24_0_I1275 (.CO(N3670), .S(N3340), .A(N3648), .B(N3117), .CI(N2574));
ADDFX1 inst_cellmath__24_0_I1276 (.CO(N2605), .S(N2262), .A(N3371), .B(N3234), .CI(N3527));
ADDFX1 inst_cellmath__24_0_I1277 (.CO(N3279), .S(N2944), .A(N3255), .B(N3313), .CI(N2782));
ADDFX1 inst_cellmath__24_0_I1278 (.CO(N2747), .S(N2309), .A(N3340), .B(N2262), .CI(N2376));
ADDFX1 inst_cellmath__24_0_I1279 (.CO(N2402), .S(N3616), .A(N2944), .B(N2522), .CI(N2309));
ADDFX1 inst_cellmath__24_0_I1280 (.CO(N3425), .S(N3084), .A(N3305), .B(N2429), .CI(N3448));
ADDFX1 inst_cellmath__24_0_I1281 (.CO(N2889), .S(N3606), .A(N3643), .B(N3504), .CI(N2225));
ADDFX1 inst_cellmath__24_0_I1282 (.CO(N2549), .S(N2202), .A(N2462), .B(N2319), .CI(N3606));
ADDFX1 inst_cellmath__24_0_I1283 (.CO(N3025), .S(N2689), .A(N2495), .B(N2363), .CI(N2817));
ADDFX1 inst_cellmath__24_0_I1284 (.CO(N2149), .S(N3365), .A(N2689), .B(N3084), .CI(N3670));
ADDFX1 inst_cellmath__24_0_I1285 (.CO(N2289), .S(N3496), .A(N2202), .B(N2605), .CI(N3279));
ADDFX1 inst_cellmath__24_0_I1286 (.CO(N2969), .S(N2630), .A(N2747), .B(N3365), .CI(N3496));
INVXL inst_cellmath__24_0_I1287 (.Y(N3158), .A(N3110));
ADDFX1 inst_cellmath__24_0_I1288 (.CO(N3640), .S(N3306), .A(N2775), .B(N2576), .CI(N3158));
ADDFX1 inst_cellmath__24_0_I1289 (.CO(N3447), .S(N3109), .A(N3039), .B(N2910), .CI(N2639));
ADDFX1 inst_cellmath__24_0_I1290 (.CO(N3580), .S(N3247), .A(N3425), .B(N3172), .CI(N2889));
ADDFX1 inst_cellmath__24_0_I1291 (.CO(N2716), .S(N2371), .A(N3109), .B(N3025), .CI(N3306));
ADDFX1 inst_cellmath__24_0_I1292 (.CO(N2174), .S(N3294), .A(N2549), .B(N3247), .CI(N2371));
ADDFX1 inst_cellmath__24_0_I1293 (.CO(N3394), .S(N3049), .A(N2149), .B(N2289), .CI(N3294));
ADDFX1 inst_cellmath__24_0_I1294 (.CO(N3189), .S(N3041), .A(N3110), .B(N2230), .CI(N3245));
ADDFX1 inst_cellmath__24_0_I1295 (.CO(N2856), .S(N2515), .A(N3449), .B(N3152), .CI(N3041));
ADDFX1 inst_cellmath__24_0_I1296 (.CO(N2656), .S(N2793), .A(N2163), .B(N3576), .CI(N2294));
ADDFX1 inst_cellmath__24_0_I1297 (.CO(N2312), .S(N3520), .A(N3447), .B(N3640), .CI(N2793));
ADDFX1 inst_cellmath__24_0_I1298 (.CO(N3663), .S(N2531), .A(N2515), .B(N3580), .CI(N2716));
ADDFX1 inst_cellmath__24_0_I1299 (.CO(N3332), .S(N2992), .A(N3520), .B(N2174), .CI(N2531));
INVXL inst_cellmath__24_0_I1300 (.Y(N3623), .A(N2914));
ADDFX1 inst_cellmath__24_0_I1301 (.CO(N2801), .S(N2456), .A(N2710), .B(N2372), .CI(N3623));
ADDFX1 inst_cellmath__24_0_I1302 (.CO(N2940), .S(N2212), .A(N2580), .B(N2847), .CI(N2974));
ADDFX1 inst_cellmath__24_0_I1303 (.CO(N2599), .S(N2256), .A(N3189), .B(N2656), .CI(N2212));
ADDFX1 inst_cellmath__24_0_I1304 (.CO(N3075), .S(N2739), .A(N2856), .B(N2456), .CI(N2312));
ADDFX1 inst_cellmath__24_0_I1305 (.CO(N2195), .S(N3418), .A(N3663), .B(N2256), .CI(N2739));
ADDFX1 inst_cellmath__24_0_I1306 (.CO(N2881), .S(N2542), .A(N2914), .B(N3581), .CI(N3050));
ADDFX1 inst_cellmath__24_0_I1307 (.CO(N2344), .S(N3503), .A(N3507), .B(N3390), .CI(N3646));
ADDFX1 inst_cellmath__24_0_I1308 (.CO(N3546), .S(N3214), .A(N2940), .B(N2801), .CI(N3503));
ADDFX1 inst_cellmath__24_0_I1309 (.CO(N2480), .S(N3687), .A(N2542), .B(N3481), .CI(N2599));
ADDFX1 inst_cellmath__24_0_I1310 (.CO(N3161), .S(N2826), .A(N3075), .B(N3214), .CI(N3687));
INVXL inst_cellmath__24_0_I1311 (.Y(N3055), .A(N2714));
ADDFX1 inst_cellmath__24_0_I1312 (.CO(N2283), .S(N3489), .A(N2642), .B(N2175), .CI(N3055));
ADDFX1 inst_cellmath__24_0_I1313 (.CO(N3634), .S(N3299), .A(N2509), .B(N2783), .CI(N2881));
ADDFX1 inst_cellmath__24_0_I1314 (.CO(N3105), .S(N3197), .A(N3489), .B(N2344), .CI(N3299));
ADDFX1 inst_cellmath__24_0_I1315 (.CO(N2767), .S(N2421), .A(N2480), .B(N3546), .CI(N3197));
ADDFX1 inst_cellmath__24_0_I1316 (.CO(N2568), .S(N2945), .A(N2714), .B(N3395), .CI(N2857));
ADDFX1 inst_cellmath__24_0_I1317 (.CO(N2224), .S(N3442), .A(N3321), .B(N2273), .CI(N2945));
ADDFX1 inst_cellmath__24_0_I1318 (.CO(N2709), .S(N2366), .A(N2283), .B(N3451), .CI(N3634));
ADDFX1 inst_cellmath__24_0_I1319 (.CO(N3386), .S(N3044), .A(N2366), .B(N3442), .CI(N3105));
INVXL inst_cellmath__24_0_I1320 (.Y(N2488), .A(N2516));
ADDFX1 inst_cellmath__24_0_I1321 (.CO(N2506), .S(N2167), .A(N2583), .B(N3518), .CI(N2488));
ADDFX1 inst_cellmath__24_0_I1322 (.CO(N3325), .S(N2983), .A(N2568), .B(N2442), .CI(N2167));
ADDFX1 inst_cellmath__24_0_I1323 (.CO(N2447), .S(N3656), .A(N2709), .B(N2224), .CI(N2983));
ADDFX1 inst_cellmath__24_0_I1324 (.CO(N3130), .S(N2797), .A(N2516), .B(N3190), .CI(N2657));
ADDFX1 inst_cellmath__24_0_I1325 (.CO(N3269), .S(N2931), .A(N2615), .B(N3256), .CI(N2797));
ADDFX1 inst_cellmath__24_0_I1326 (.CO(N2389), .S(N3601), .A(N2931), .B(N2506), .CI(N3325));
INVXL inst_cellmath__24_0_I1327 (.Y(N2430), .A(N2313));
ADDFX1 inst_cellmath__24_0_I1328 (.CO(N3068), .S(N2732), .A(N2377), .B(N3333), .CI(N2430));
ADDFX1 inst_cellmath__24_0_I1329 (.CO(N2875), .S(N2536), .A(N2732), .B(N3130), .CI(N3269));
ADDFX1 inst_cellmath__24_0_I1330 (.CO(N3011), .S(N2676), .A(N2313), .B(N2990), .CI(N2454));
ADDFX1 inst_cellmath__24_0_I1331 (.CO(N3679), .S(N3352), .A(N2676), .B(N2955), .CI(N3068));
ADDFX1 inst_cellmath__24_0_I1332 (.CO(N2614), .S(N2275), .A(N3134), .B(N3136), .CI(N3011));
XNOR2X1 inst_cellmath__24_0_I1333 (.Y(N2761), .A(N2938), .B(N3134));
AND2XL inst_cellmath__24_0_I1334 (.Y(N3435), .A(b_man[1]), .B(N2292));
NOR2XL inst_cellmath__24_0_I1335 (.Y(N2560), .A(N2231), .B(N3290));
NAND2XL inst_cellmath__24_0_I1336 (.Y(N2898), .A(N2231), .B(N3290));
NOR2XL inst_cellmath__24_0_I1337 (.Y(N3232), .A(N3626), .B(N2412));
NAND2XL inst_cellmath__24_0_I1338 (.Y(N3568), .A(N3626), .B(N2412));
NOR2XL inst_cellmath__24_0_I1339 (.Y(N2361), .A(N3095), .B(N2215));
NAND2XL inst_cellmath__24_0_I1340 (.Y(N2702), .A(N3095), .B(N2215));
NOR2XL inst_cellmath__24_0_I1341 (.Y(N3036), .A(N2561), .B(N3569));
NAND2XL inst_cellmath__24_0_I1342 (.Y(N3376), .A(N2561), .B(N3569));
NOR2XL inst_cellmath__24_0_I1343 (.Y(N2162), .A(N2362), .B(N3377));
NAND2XL inst_cellmath__24_0_I1344 (.Y(N2498), .A(N2362), .B(N3377));
NOR2XL inst_cellmath__24_0_I1345 (.Y(N2845), .A(N2161), .B(N3649));
NAND2XL inst_cellmath__24_0_I1346 (.Y(N3176), .A(N2161), .B(N3649));
NOR2XL inst_cellmath__24_0_I1347 (.Y(N3505), .A(N2439), .B(N2588));
NAND2XL inst_cellmath__24_0_I1348 (.Y(N2298), .A(N2439), .B(N2588));
NOR2XL inst_cellmath__24_0_I1349 (.Y(N2640), .A(N2926), .B(N3531));
NAND2XL inst_cellmath__24_0_I1350 (.Y(N2976), .A(N2926), .B(N3531));
NOR2XL inst_cellmath__24_0_I1351 (.Y(N3318), .A(N2327), .B(N2948));
NAND2XL inst_cellmath__24_0_I1352 (.Y(N3651), .A(N2327), .B(N2948));
NOR2XL inst_cellmath__24_0_I1353 (.Y(N2438), .A(N3283), .B(N2355));
NAND2XL inst_cellmath__24_0_I1354 (.Y(N2787), .A(N3283), .B(N2355));
NOR2XL inst_cellmath__24_0_I1355 (.Y(N3123), .A(N2694), .B(N2433));
NAND2XL inst_cellmath__24_0_I1356 (.Y(N3455), .A(N2694), .B(N2433));
NOR2XL inst_cellmath__24_0_I1357 (.Y(N2244), .A(N2780), .B(N2317));
NAND2XL inst_cellmath__24_0_I1358 (.Y(N2590), .A(N2780), .B(N2317));
NOR2XL inst_cellmath__24_0_I1359 (.Y(N2925), .A(N2663), .B(N2744));
NAND2XL inst_cellmath__24_0_I1360 (.Y(N3262), .A(N2663), .B(N2744));
NOR2XL inst_cellmath__24_0_I1361 (.Y(N3594), .A(N3082), .B(N3165));
NAND2XL inst_cellmath__24_0_I1362 (.Y(N2381), .A(N3082), .B(N3165));
NOR2X1 inst_cellmath__24_0_I1363 (.Y(N2726), .A(N3494), .B(N2513));
NAND2XL inst_cellmath__24_0_I1364 (.Y(N3063), .A(N3494), .B(N2513));
NOR2XL inst_cellmath__24_0_I1365 (.Y(N3405), .A(N2854), .B(N3415));
NAND2XL inst_cellmath__24_0_I1366 (.Y(N2186), .A(N2854), .B(N3415));
NOR2XL inst_cellmath__24_0_I1367 (.Y(N2527), .A(N2193), .B(N2960));
NAND2XL inst_cellmath__24_0_I1368 (.Y(N2867), .A(N2193), .B(N2960));
AND2XL inst_cellmath__24_0_I1369 (.Y(N2326), .A(N2217), .B(N3435));
INVXL inst_cellmath__24_0_I1370 (.Y(N2423), .A(N2560));
INVXL inst_cellmath__24_0_I1371 (.Y(N2769), .A(N2898));
OAI21XL inst_cellmath__24_0_I1372 (.Y(N2607), .A0(N2769), .A1(N2326), .B0(N2423));
AOI21XL inst_cellmath__24_0_I1373 (.Y(N2208), .A0(N3568), .A1(N2607), .B0(N3232));
INVXL inst_cellmath__24_0_I1374 (.Y(N3241), .A(N2361));
INVXL inst_cellmath__24_0_I1375 (.Y(N3574), .A(N2702));
OAI21XL inst_cellmath__24_0_I1376 (.Y(N3170), .A0(N3574), .A1(N2208), .B0(N3241));
AOI21XL inst_cellmath__24_0_I1377 (.Y(N2582), .A0(N3376), .A1(N3170), .B0(N3036));
INVXL inst_cellmath__24_0_I1378 (.Y(N2307), .A(N2162));
INVXL inst_cellmath__24_0_I1379 (.Y(N2650), .A(N2498));
OAI21XL inst_cellmath__24_0_I1380 (.Y(N3337), .A0(N2650), .A1(N2582), .B0(N2307));
AO21XL inst_cellmath__24_0_I1381 (.Y(N3270), .A0(N2298), .A1(N2845), .B0(N3505));
AOI21XL inst_cellmath__24_0_I1382 (.Y(N2147), .A0(N3176), .A1(N3337), .B0(N2845));
AOI31X1 inst_cellmath__24_0_I1383 (.Y(N2834), .A0(N2298), .A1(N3176), .A2(N3337), .B0(N3270));
INVXL inst_cellmath__24_0_I1384 (.Y(N3208), .A(N2640));
INVXL inst_cellmath__24_0_I1385 (.Y(N3539), .A(N2976));
OAI21XL inst_cellmath__24_0_I1386 (.Y(N2514), .A0(N3539), .A1(N2834), .B0(N3208));
AO21XL inst_cellmath__24_0_I1387 (.Y(N3628), .A0(N2787), .A1(N3318), .B0(N2438));
AND2XL inst_cellmath__24_0_I1388 (.Y(N2414), .A(N2787), .B(N3651));
AOI21XL inst_cellmath__24_0_I1389 (.Y(N3360), .A0(N3651), .A1(N2514), .B0(N3318));
AOI21X1 inst_cellmath__24_0_I1390 (.Y(N2478), .A0(N2414), .A1(N2514), .B0(N3628));
AOI21XL inst_cellmath__24_0_I1392 (.Y(N2281), .A0(N2590), .A1(N3123), .B0(N2244));
NAND2XL inst_cellmath__24_0_I1393 (.Y(N2621), .A(N2590), .B(N3455));
OAI21X1 inst_cellmath__24_0_I1394 (.Y(N2445), .A0(N2621), .A1(N2478), .B0(N2281));
AO21XL inst_cellmath__24_0_I1395 (.Y(N2928), .A0(N2381), .A1(N2925), .B0(N3594));
AND2XL inst_cellmath__24_0_I1396 (.Y(N3264), .A(N2381), .B(N3262));
NOR2BX1 inst_cellmath__24_0_I3658 (.Y(N3560), .AN(N3455), .B(N2478));
NOR2XL inst_cellmath__24_0_I1398 (.Y(N3006), .A(N3560), .B(N3123));
AOI21XL inst_cellmath__24_0_I1399 (.Y(N2895), .A0(N3262), .A1(N2445), .B0(N2925));
AOI21X1 inst_cellmath__24_0_I1400 (.Y(N3565), .A0(N3264), .A1(N2445), .B0(N2928));
AOI21XL inst_cellmath__24_0_I1401 (.Y(N3374), .A0(N2186), .A1(N2726), .B0(N3405));
NAND2XL inst_cellmath__24_0_I1402 (.Y(N2160), .A(N2186), .B(N3063));
INVXL inst_cellmath__24_0_I1403 (.Y(N3148), .A(N2867));
INVXL inst_cellmath__24_0_I1404 (.Y(N3285), .A(N2726));
INVXL inst_cellmath__24_0_I1405 (.Y(N3621), .A(N3063));
NOR2XL inst_cellmath__24_0_I1406 (.Y(N2842), .A(N3148), .B(N3374));
NOR2XL inst_cellmath__24_0_I1407 (.Y(N3091), .A(N2842), .B(N2527));
OAI21XL inst_cellmath__24_0_I1408 (.Y(N2552), .A0(N3621), .A1(N3565), .B0(N3285));
OAI21XL inst_cellmath__24_0_I1409 (.Y(N3224), .A0(N2160), .A1(N3565), .B0(N3374));
OAI31X1 inst_cellmath__24_0_I1410 (.Y(N3388), .A0(N3148), .A1(N2160), .A2(N3565), .B0(N3091));
NAND2BXL inst_cellmath__24_0_I1411 (.Y(N3308), .AN(N2560), .B(N2898));
NAND2BXL inst_cellmath__24_0_I1412 (.Y(N2777), .AN(N3232), .B(N3568));
NAND2BXL inst_cellmath__24_0_I1413 (.Y(N2233), .AN(N2361), .B(N2702));
NAND2BXL inst_cellmath__24_0_I1414 (.Y(N3248), .AN(N3036), .B(N3376));
NAND2BXL inst_cellmath__24_0_I1415 (.Y(N2717), .AN(N2162), .B(N2498));
NAND2BXL inst_cellmath__24_0_I1416 (.Y(N2177), .AN(N2845), .B(N3176));
NAND2BXL inst_cellmath__24_0_I1417 (.Y(N3191), .AN(N3505), .B(N2298));
NAND2BXL inst_cellmath__24_0_I1418 (.Y(N2660), .AN(N2640), .B(N2976));
NAND2BXL inst_cellmath__24_0_I1419 (.Y(N3666), .AN(N3318), .B(N3651));
NAND2BXL inst_cellmath__24_0_I1420 (.Y(N3138), .AN(N2438), .B(N2787));
NAND2BXL inst_cellmath__24_0_I1421 (.Y(N2601), .AN(N3123), .B(N3455));
NAND2BXL inst_cellmath__24_0_I1422 (.Y(N3610), .AN(N2244), .B(N2590));
NAND2BXL inst_cellmath__24_0_I1423 (.Y(N3077), .AN(N2925), .B(N3262));
NAND2BXL inst_cellmath__24_0_I1424 (.Y(N2543), .AN(N3594), .B(N2381));
NAND2BXL inst_cellmath__24_0_I1425 (.Y(N3548), .AN(N2726), .B(N3063));
NAND2BXL inst_cellmath__24_0_I1426 (.Y(N3020), .AN(N3405), .B(N2186));
NAND2BXL inst_cellmath__24_0_I1427 (.Y(N2481), .AN(N2527), .B(N2867));
XOR2XL inst_cellmath__24_0_I1428 (.Y(inst_cellmath__24[0]), .A(b_man[1]), .B(N2292));
XOR2XL inst_cellmath__24_0_I1429 (.Y(inst_cellmath__24[1]), .A(N3435), .B(N2217));
XNOR2X1 inst_cellmath__24_0_I1430 (.Y(inst_cellmath__24[2]), .A(N2326), .B(N3308));
XOR2XL inst_cellmath__24_0_I1431 (.Y(inst_cellmath__24[3]), .A(N2607), .B(N2777));
XNOR2X1 inst_cellmath__24_0_I1432 (.Y(inst_cellmath__24[4]), .A(N2208), .B(N2233));
XOR2XL inst_cellmath__24_0_I1433 (.Y(inst_cellmath__24[5]), .A(N3170), .B(N3248));
XNOR2X1 inst_cellmath__24_0_I1434 (.Y(inst_cellmath__24[6]), .A(N2582), .B(N2717));
XOR2XL inst_cellmath__24_0_I1435 (.Y(inst_cellmath__24[7]), .A(N3337), .B(N2177));
XNOR2X1 inst_cellmath__24_0_I1436 (.Y(inst_cellmath__24[8]), .A(N2147), .B(N3191));
XNOR2X1 inst_cellmath__24_0_I1437 (.Y(inst_cellmath__24[9]), .A(N2834), .B(N2660));
XOR2XL inst_cellmath__24_0_I1438 (.Y(inst_cellmath__24[10]), .A(N2514), .B(N3666));
XNOR2X1 inst_cellmath__24_0_I1439 (.Y(inst_cellmath__24[11]), .A(N3360), .B(N3138));
XNOR2X1 inst_cellmath__24_0_I1440 (.Y(inst_cellmath__24[12]), .A(N2478), .B(N2601));
XNOR2X1 inst_cellmath__24_0_I1441 (.Y(inst_cellmath__24[13]), .A(N3006), .B(N3610));
XOR2XL inst_cellmath__24_0_I1442 (.Y(inst_cellmath__24[14]), .A(N2445), .B(N3077));
XNOR2X1 inst_cellmath__24_0_I1443 (.Y(inst_cellmath__24[15]), .A(N2895), .B(N2543));
XNOR2X1 inst_cellmath__24_0_I1444 (.Y(inst_cellmath__24[16]), .A(N3565), .B(N3548));
XOR2XL inst_cellmath__24_0_I1445 (.Y(inst_cellmath__24[17]), .A(N2552), .B(N3020));
XOR2XL inst_cellmath__24_0_I1446 (.Y(inst_cellmath__24[18]), .A(N3224), .B(N2481));
OR2XL inst_cellmath__24_0_I1447 (.Y(N2578), .A(N3296), .B(N2849));
XOR2XL inst_cellmath__24_0_I1448 (.Y(N2851), .A(N3296), .B(N2849));
OR2XL inst_cellmath__24_0_I1449 (.Y(N3397), .A(N3182), .B(N3409));
XOR2XL inst_cellmath__24_0_I1450 (.Y(N3512), .A(N3182), .B(N3409));
XOR2XL inst_cellmath__24_0_I1451 (.Y(N2651), .A(N2188), .B(N2558));
XOR2XL inst_cellmath__24_0_I1452 (.Y(N3327), .A(N2896), .B(N2922));
OR2XL inst_cellmath__24_0_I1453 (.Y(N2741), .A(N3259), .B(N2404));
XOR2XL inst_cellmath__24_0_I1454 (.Y(N2451), .A(N3259), .B(N2404));
OR2XL inst_cellmath__24_0_I1455 (.Y(N3547), .A(N2750), .B(N3309));
XOR2XL inst_cellmath__24_0_I1456 (.Y(N3131), .A(N2750), .B(N3309));
OR2XL inst_cellmath__24_0_I1457 (.Y(N2827), .A(N3642), .B(N3139));
XOR2XL inst_cellmath__24_0_I1458 (.Y(N2251), .A(N3642), .B(N3139));
OR2XL inst_cellmath__24_0_I1459 (.Y(N3635), .A(N3467), .B(N3163));
XOR2XL inst_cellmath__24_0_I1460 (.Y(N2934), .A(N3467), .B(N3163));
OR2XL inst_cellmath__24_0_I1461 (.Y(N2908), .A(N3491), .B(N2508));
XOR2XL inst_cellmath__24_0_I1462 (.Y(N3604), .A(N3491), .B(N2508));
OR2XL inst_cellmath__24_0_I1463 (.Y(N2168), .A(N2852), .B(N3540));
XOR2XL inst_cellmath__24_0_I1464 (.Y(N2734), .A(N2852), .B(N3540));
OR2XL inst_cellmath__24_0_I1465 (.Y(N2985), .A(N2337), .B(N3437));
XOR2XL inst_cellmath__24_0_I1466 (.Y(N3414), .A(N2337), .B(N3437));
OR2XL inst_cellmath__24_0_I1467 (.Y(N2250), .A(N2220), .B(N2384));
XOR2XL inst_cellmath__24_0_I1468 (.Y(N2538), .A(N2220), .B(N2384));
OR2XL inst_cellmath__24_0_I1469 (.Y(N3069), .A(N2729), .B(N3477));
XOR2XL inst_cellmath__24_0_I1470 (.Y(N3209), .A(N2729), .B(N3477));
OR2XL inst_cellmath__24_0_I1471 (.Y(N2336), .A(N2269), .B(N2293));
XOR2XL inst_cellmath__24_0_I1472 (.Y(N2339), .A(N2269), .B(N2293));
OR2XL inst_cellmath__24_0_I1473 (.Y(N3154), .A(N2637), .B(N2862));
XOR2XL inst_cellmath__24_0_I1474 (.Y(N3014), .A(N2637), .B(N2862));
OR2XL inst_cellmath__24_0_I1475 (.Y(N2413), .A(N3196), .B(N3616));
XOR2XL inst_cellmath__24_0_I1476 (.Y(N3682), .A(N3196), .B(N3616));
OR2XL inst_cellmath__24_0_I1477 (.Y(N3233), .A(N2402), .B(N2630));
XOR2XL inst_cellmath__24_0_I1478 (.Y(N2821), .A(N2402), .B(N2630));
OR2XL inst_cellmath__24_0_I1479 (.Y(N2501), .A(N2969), .B(N3049));
XOR2XL inst_cellmath__24_0_I1480 (.Y(N3483), .A(N2969), .B(N3049));
OR2XL inst_cellmath__24_0_I1481 (.Y(N3320), .A(N3394), .B(N2992));
XOR2XL inst_cellmath__24_0_I1482 (.Y(N2617), .A(N3394), .B(N2992));
OR2XL inst_cellmath__24_0_I1483 (.Y(N2591), .A(N3332), .B(N3418));
XOR2XL inst_cellmath__24_0_I1484 (.Y(N3293), .A(N3332), .B(N3418));
OR2XL inst_cellmath__24_0_I1485 (.Y(N3407), .A(N2195), .B(N2826));
XOR2XL inst_cellmath__24_0_I1486 (.Y(N2415), .A(N2195), .B(N2826));
OR2XL inst_cellmath__24_0_I1487 (.Y(N2672), .A(N3161), .B(N2421));
XOR2XL inst_cellmath__24_0_I1488 (.Y(N3100), .A(N3161), .B(N2421));
OR2XL inst_cellmath__24_0_I1489 (.Y(N3475), .A(N3044), .B(N2767));
XOR2XL inst_cellmath__24_0_I1490 (.Y(N2219), .A(N3044), .B(N2767));
OR2XL inst_cellmath__24_0_I1491 (.Y(N2755), .A(N3386), .B(N3656));
XOR2XL inst_cellmath__24_0_I1492 (.Y(N2900), .A(N3386), .B(N3656));
OR2XL inst_cellmath__24_0_I1493 (.Y(N3561), .A(N2447), .B(N3601));
XOR2XL inst_cellmath__24_0_I1494 (.Y(N3571), .A(N2447), .B(N3601));
OR2XL inst_cellmath__24_0_I1495 (.Y(N2840), .A(N2536), .B(N2389));
XOR2XL inst_cellmath__24_0_I1496 (.Y(N2704), .A(N2536), .B(N2389));
OR2XL inst_cellmath__24_0_I1497 (.Y(N3645), .A(N3352), .B(N2875));
XOR2XL inst_cellmath__24_0_I1498 (.Y(N3379), .A(N3352), .B(N2875));
OR2XL inst_cellmath__24_0_I1499 (.Y(N2917), .A(N2275), .B(N3679));
XOR2XL inst_cellmath__24_0_I1500 (.Y(N2503), .A(N2275), .B(N3679));
XNOR2X1 inst_cellmath__24_0_I1501 (.Y(N3178), .A(N2614), .B(N2761));
OAI2BB1X1 inst_cellmath__24_0_I1502 (.Y(N2643), .A0N(N2851), .A1N(N3388), .B0(N2578));
OAI2BB1X1 inst_cellmath__24_0_I1503 (.Y(N3124), .A0N(N3512), .A1N(N2643), .B0(N3397));
OAI2BB2XL inst_cellmath__24_0_I1504 (.Y(N2728), .A0N(N2651), .A1N(N3124), .B0(N2188), .B1(N2558));
OAI2BB2XL inst_cellmath__24_0_I1505 (.Y(N3007), .A0N(N3327), .A1N(N2728), .B0(N2896), .B1(N2922));
OAI2BB1X1 inst_cellmath__24_0_I1506 (.Y(N2409), .A0N(N2451), .A1N(N3007), .B0(N2741));
OAI2BB1X1 inst_cellmath__24_0_I1507 (.Y(N2494), .A0N(N3131), .A1N(N2409), .B0(N3547));
OAI2BB1X1 inst_cellmath__24_0_I1508 (.Y(N3254), .A0N(N2251), .A1N(N2494), .B0(N2827));
OAI2BB1X1 inst_cellmath__24_0_I1509 (.Y(N3144), .A0N(N2934), .A1N(N3254), .B0(N3635));
OAI2BB1X1 inst_cellmath__24_0_I1510 (.Y(N2151), .A0N(N3604), .A1N(N3144), .B0(N2908));
OAI2BB1X1 inst_cellmath__24_0_I1511 (.Y(N3393), .A0N(N2734), .A1N(N2151), .B0(N2168));
OAI2BB1X1 inst_cellmath__24_0_I1512 (.Y(N2197), .A0N(N3414), .A1N(N3393), .B0(N2985));
OAI2BB1X1 inst_cellmath__24_0_I1513 (.Y(N3239), .A0N(N2538), .A1N(N2197), .B0(N2250));
OAI2BB1X1 inst_cellmath__24_0_I1514 (.Y(N3412), .A0N(N3209), .A1N(N3239), .B0(N3069));
OAI2BB1X1 inst_cellmath__24_0_I1515 (.Y(N2701), .A0N(N2339), .A1N(N3412), .B0(N2336));
OAI2BB1X1 inst_cellmath__24_0_I1516 (.Y(N2670), .A0N(N3014), .A1N(N2701), .B0(N3154));
OAI2BB1X1 inst_cellmath__24_0_I1517 (.Y(N3310), .A0N(N3682), .A1N(N2670), .B0(N2413));
OAI2BB1X1 inst_cellmath__24_0_I1518 (.Y(N3081), .A0N(N2821), .A1N(N3310), .B0(N3233));
OAI2BB1X1 inst_cellmath__24_0_I1519 (.Y(N3516), .A0N(N3483), .A1N(N3081), .B0(N2501));
OAI2BB1X1 inst_cellmath__24_0_I1520 (.Y(N3104), .A0N(N2617), .A1N(N3516), .B0(N3320));
OAI2BB1X1 inst_cellmath__24_0_I1521 (.Y(N3349), .A0N(N3293), .A1N(N3104), .B0(N2591));
OAI2BB1X1 inst_cellmath__24_0_I1522 (.Y(N2723), .A0N(N2415), .A1N(N3349), .B0(N3407));
OAI2BB1X1 inst_cellmath__24_0_I1523 (.Y(N2776), .A0N(N3100), .A1N(N2723), .B0(N2672));
OAI2BB1X1 inst_cellmath__24_0_I1524 (.Y(N3493), .A0N(N2219), .A1N(N2776), .B0(N3475));
OAI2BB1X1 inst_cellmath__24_0_I1525 (.Y(N3356), .A0N(N2900), .A1N(N3493), .B0(N2755));
OAI2BB1X1 inst_cellmath__24_0_I1526 (.Y(N2331), .A0N(N3571), .A1N(N3356), .B0(N3561));
OAI2BB1X1 inst_cellmath__24_0_I1527 (.Y(N3526), .A0N(N2704), .A1N(N2331), .B0(N2840));
OAI2BB1X1 inst_cellmath__24_0_I1528 (.Y(N2315), .A0N(N3379), .A1N(N3526), .B0(N3645));
OAI2BB1X1 inst_cellmath__24_0_I1529 (.Y(N3326), .A0N(N2503), .A1N(N2315), .B0(N2917));
XNOR2X1 inst_cellmath__24_0_I1530 (.Y(inst_cellmath__24[19]), .A(N3388), .B(N2851));
XNOR2X1 inst_cellmath__24_0_I1531 (.Y(inst_cellmath__24[20]), .A(N2643), .B(N3512));
XNOR2X1 inst_cellmath__24_0_I1532 (.Y(inst_cellmath__24[21]), .A(N3124), .B(N2651));
XNOR2X1 inst_cellmath__24_0_I1533 (.Y(inst_cellmath__24[22]), .A(N2728), .B(N3327));
XNOR2X1 inst_cellmath__24_0_I1534 (.Y(inst_cellmath__24[23]), .A(N3007), .B(N2451));
XNOR2X1 inst_cellmath__24_0_I1535 (.Y(inst_cellmath__24[24]), .A(N2409), .B(N3131));
XNOR2X1 inst_cellmath__24_0_I1536 (.Y(inst_cellmath__24[25]), .A(N2494), .B(N2251));
XNOR2X1 inst_cellmath__24_0_I1537 (.Y(inst_cellmath__24[26]), .A(N3254), .B(N2934));
XNOR2X1 inst_cellmath__24_0_I1538 (.Y(inst_cellmath__24[27]), .A(N3144), .B(N3604));
XNOR2X1 inst_cellmath__24_0_I1539 (.Y(inst_cellmath__24[28]), .A(N2151), .B(N2734));
XNOR2X1 inst_cellmath__24_0_I1540 (.Y(inst_cellmath__24[29]), .A(N3393), .B(N3414));
XNOR2X1 inst_cellmath__24_0_I1541 (.Y(inst_cellmath__24[30]), .A(N2197), .B(N2538));
XNOR2X1 inst_cellmath__24_0_I1542 (.Y(inst_cellmath__24[31]), .A(N3239), .B(N3209));
XNOR2X1 inst_cellmath__24_0_I1543 (.Y(inst_cellmath__24[32]), .A(N3412), .B(N2339));
XNOR2X1 inst_cellmath__24_0_I1544 (.Y(inst_cellmath__24[33]), .A(N2701), .B(N3014));
XNOR2X1 inst_cellmath__24_0_I1545 (.Y(inst_cellmath__24[34]), .A(N2670), .B(N3682));
XNOR2X1 inst_cellmath__24_0_I1546 (.Y(inst_cellmath__24[35]), .A(N3310), .B(N2821));
XNOR2X1 inst_cellmath__24_0_I1547 (.Y(inst_cellmath__24[36]), .A(N3081), .B(N3483));
XNOR2X1 inst_cellmath__24_0_I1548 (.Y(inst_cellmath__24[37]), .A(N3516), .B(N2617));
XNOR2X1 inst_cellmath__24_0_I1549 (.Y(inst_cellmath__24[38]), .A(N3104), .B(N3293));
XNOR2X1 inst_cellmath__24_0_I1550 (.Y(inst_cellmath__24[39]), .A(N3349), .B(N2415));
XNOR2X1 inst_cellmath__24_0_I1551 (.Y(inst_cellmath__24[40]), .A(N2723), .B(N3100));
XNOR2X1 inst_cellmath__24_0_I1552 (.Y(inst_cellmath__24[41]), .A(N2776), .B(N2219));
XNOR2X1 inst_cellmath__24_0_I1553 (.Y(inst_cellmath__24[42]), .A(N3493), .B(N2900));
XNOR2X1 inst_cellmath__24_0_I1554 (.Y(inst_cellmath__24[43]), .A(N3356), .B(N3571));
XNOR2X1 inst_cellmath__24_0_I1555 (.Y(inst_cellmath__24[44]), .A(N2331), .B(N2704));
XNOR2X1 inst_cellmath__24_0_I1556 (.Y(inst_cellmath__24[45]), .A(N3526), .B(N3379));
XNOR2X1 inst_cellmath__24_0_I1557 (.Y(inst_cellmath__24[46]), .A(N2315), .B(N2503));
XOR2XL inst_cellmath__24_0_I1558 (.Y(inst_cellmath__24[47]), .A(N3326), .B(N3178));
BUFX2 inst_cellmath__25_0_I1559 (.Y(N5224), .A(inst_cellmath__24[47]));
INVX2 inst_cellmath__25_0_I3631 (.Y(N8368), .A(N5224));
INVX2 inst_cellmath__25_0_I3639 (.Y(N8376), .A(N8368));
INVX2 inst_cellmath__25_0_I3636 (.Y(N8373), .A(N8368));
AND2XL inst_cellmath__25_0_I1560 (.Y(inst_cellmath__25[0]), .A(N8376), .B(inst_cellmath__24[0]));
MX2XL inst_cellmath__25_0_I1561 (.Y(inst_cellmath__25[1]), .A(inst_cellmath__24[0]), .B(inst_cellmath__24[1]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1562 (.Y(inst_cellmath__25[2]), .A(inst_cellmath__24[1]), .B(inst_cellmath__24[2]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1563 (.Y(inst_cellmath__25[3]), .A(inst_cellmath__24[2]), .B(inst_cellmath__24[3]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1564 (.Y(inst_cellmath__25[4]), .A(inst_cellmath__24[3]), .B(inst_cellmath__24[4]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1565 (.Y(inst_cellmath__25[5]), .A(inst_cellmath__24[4]), .B(inst_cellmath__24[5]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1566 (.Y(inst_cellmath__25[6]), .A(inst_cellmath__24[5]), .B(inst_cellmath__24[6]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1567 (.Y(inst_cellmath__25[7]), .A(inst_cellmath__24[6]), .B(inst_cellmath__24[7]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1568 (.Y(inst_cellmath__25[8]), .A(inst_cellmath__24[7]), .B(inst_cellmath__24[8]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1569 (.Y(inst_cellmath__25[9]), .A(inst_cellmath__24[8]), .B(inst_cellmath__24[9]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1570 (.Y(inst_cellmath__25[10]), .A(inst_cellmath__24[9]), .B(inst_cellmath__24[10]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1571 (.Y(inst_cellmath__25[11]), .A(inst_cellmath__24[10]), .B(inst_cellmath__24[11]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1572 (.Y(inst_cellmath__25[12]), .A(inst_cellmath__24[11]), .B(inst_cellmath__24[12]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1573 (.Y(inst_cellmath__25[13]), .A(inst_cellmath__24[12]), .B(inst_cellmath__24[13]), .S0(N5224));
MX2XL inst_cellmath__25_0_I1574 (.Y(inst_cellmath__25[14]), .A(inst_cellmath__24[13]), .B(inst_cellmath__24[14]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1575 (.Y(inst_cellmath__25[15]), .A(inst_cellmath__24[14]), .B(inst_cellmath__24[15]), .S0(N5224));
MX2XL inst_cellmath__25_0_I1576 (.Y(inst_cellmath__25[16]), .A(inst_cellmath__24[15]), .B(inst_cellmath__24[16]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1577 (.Y(inst_cellmath__25[17]), .A(inst_cellmath__24[16]), .B(inst_cellmath__24[17]), .S0(N5224));
MX2XL inst_cellmath__25_0_I1578 (.Y(inst_cellmath__25[18]), .A(inst_cellmath__24[17]), .B(inst_cellmath__24[18]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1579 (.Y(inst_cellmath__25[19]), .A(inst_cellmath__24[18]), .B(inst_cellmath__24[19]), .S0(N5224));
MX2XL inst_cellmath__25_0_I1580 (.Y(inst_cellmath__25[20]), .A(inst_cellmath__24[19]), .B(inst_cellmath__24[20]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1581 (.Y(inst_cellmath__25[21]), .A(inst_cellmath__24[20]), .B(inst_cellmath__24[21]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1582 (.Y(inst_cellmath__25[22]), .A(inst_cellmath__24[21]), .B(inst_cellmath__24[22]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1583 (.Y(inst_cellmath__25[23]), .A(inst_cellmath__24[22]), .B(inst_cellmath__24[23]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1584 (.Y(inst_cellmath__25[24]), .A(inst_cellmath__24[23]), .B(inst_cellmath__24[24]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1585 (.Y(inst_cellmath__25[25]), .A(inst_cellmath__24[24]), .B(inst_cellmath__24[25]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1586 (.Y(inst_cellmath__25[26]), .A(inst_cellmath__24[25]), .B(inst_cellmath__24[26]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1587 (.Y(inst_cellmath__25[27]), .A(inst_cellmath__24[26]), .B(inst_cellmath__24[27]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1588 (.Y(inst_cellmath__25[28]), .A(inst_cellmath__24[27]), .B(inst_cellmath__24[28]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1589 (.Y(inst_cellmath__25[29]), .A(inst_cellmath__24[28]), .B(inst_cellmath__24[29]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1590 (.Y(inst_cellmath__25[30]), .A(inst_cellmath__24[29]), .B(inst_cellmath__24[30]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1591 (.Y(inst_cellmath__25[31]), .A(inst_cellmath__24[30]), .B(inst_cellmath__24[31]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1592 (.Y(inst_cellmath__25[32]), .A(inst_cellmath__24[31]), .B(inst_cellmath__24[32]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1593 (.Y(inst_cellmath__25[33]), .A(inst_cellmath__24[32]), .B(inst_cellmath__24[33]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1594 (.Y(inst_cellmath__25[34]), .A(inst_cellmath__24[33]), .B(inst_cellmath__24[34]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1595 (.Y(inst_cellmath__25[35]), .A(inst_cellmath__24[34]), .B(inst_cellmath__24[35]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1596 (.Y(inst_cellmath__25[36]), .A(inst_cellmath__24[35]), .B(inst_cellmath__24[36]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1597 (.Y(inst_cellmath__25[37]), .A(inst_cellmath__24[36]), .B(inst_cellmath__24[37]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1598 (.Y(inst_cellmath__25[38]), .A(inst_cellmath__24[37]), .B(inst_cellmath__24[38]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1599 (.Y(inst_cellmath__25[39]), .A(inst_cellmath__24[38]), .B(inst_cellmath__24[39]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1600 (.Y(inst_cellmath__25[40]), .A(inst_cellmath__24[39]), .B(inst_cellmath__24[40]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1601 (.Y(inst_cellmath__25[41]), .A(inst_cellmath__24[40]), .B(inst_cellmath__24[41]), .S0(N8373));
MX2XL inst_cellmath__25_0_I1602 (.Y(inst_cellmath__25[42]), .A(inst_cellmath__24[41]), .B(inst_cellmath__24[42]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1603 (.Y(inst_cellmath__25[43]), .A(inst_cellmath__24[42]), .B(inst_cellmath__24[43]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1604 (.Y(inst_cellmath__25[44]), .A(inst_cellmath__24[43]), .B(inst_cellmath__24[44]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1605 (.Y(inst_cellmath__25[45]), .A(inst_cellmath__24[44]), .B(inst_cellmath__24[45]), .S0(N8376));
MX2XL inst_cellmath__25_0_I1606 (.Y(inst_cellmath__25[46]), .A(inst_cellmath__24[45]), .B(inst_cellmath__24[46]), .S0(N8376));
NOR2XL inst_cellmath__25_0_I1607 (.Y(inst_cellmath__25[47]), .A(N8376), .B(inst_cellmath__24[46]));
INVXL inst_cellmath__45_0_I1608 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__25[24]));
NAND2XL inst_cellmath__45_0_I1609 (.Y(N5411), .A(inst_cellmath__25[26]), .B(inst_cellmath__25[25]));
NOR2XL inst_cellmath__45_0_I1610 (.Y(N5387), .A(N5411), .B(inst_cellmath__45[0]));
NAND2XL inst_cellmath__45_0_I1611 (.Y(N5416), .A(inst_cellmath__25[28]), .B(inst_cellmath__25[27]));
NAND2XL inst_cellmath__45_0_I1612 (.Y(N5405), .A(inst_cellmath__25[30]), .B(inst_cellmath__25[29]));
NOR2XL inst_cellmath__45_0_I1613 (.Y(N5378), .A(N5405), .B(N5416));
NAND2XL inst_cellmath__45_0_I1614 (.Y(N5375), .A(inst_cellmath__25[27]), .B(N5387));
NAND2BXL inst_cellmath__45_0_I1615 (.Y(N5346), .AN(N5416), .B(N5387));
NAND3BXL inst_cellmath__45_0_I1616 (.Y(N5406), .AN(N5416), .B(inst_cellmath__25[29]), .C(N5387));
NAND2X1 inst_cellmath__45_0_I1617 (.Y(N5373), .A(N5378), .B(N5387));
NAND2XL inst_cellmath__45_0_I1618 (.Y(N5403), .A(inst_cellmath__25[32]), .B(inst_cellmath__25[31]));
NAND2XL inst_cellmath__45_0_I1619 (.Y(N5390), .A(inst_cellmath__25[34]), .B(inst_cellmath__25[33]));
NOR2XL inst_cellmath__45_0_I1620 (.Y(N5365), .A(N5390), .B(N5403));
NAND2XL inst_cellmath__45_0_I1621 (.Y(N5353), .A(inst_cellmath__25[36]), .B(inst_cellmath__25[35]));
NAND2XL inst_cellmath__45_0_I1622 (.Y(N5345), .A(inst_cellmath__25[38]), .B(inst_cellmath__25[37]));
NOR2XL inst_cellmath__45_0_I1623 (.Y(N5412), .A(N5345), .B(N5353));
NAND3BXL inst_cellmath__45_0_I1624 (.Y(N5419), .AN(N5353), .B(inst_cellmath__25[37]), .C(N5365));
NOR3BXL inst_cellmath__45_0_I1626 (.Y(N5363), .AN(inst_cellmath__25[33]), .B(N5403), .C(N5373));
NOR3BXL inst_cellmath__45_0_I1627 (.Y(N5359), .AN(N5365), .B(N5353), .C(N5373));
NAND2XL hyperpropagate_3_1_A_I3710 (.Y(N8402), .A(N5412), .B(N5365));
NOR2XL hyperpropagate_3_1_A_I3711 (.Y(N5392), .A(N5373), .B(N8402));
NAND2XL inst_cellmath__45_0_I1629 (.Y(N5422), .A(inst_cellmath__25[40]), .B(inst_cellmath__25[39]));
NAND2XL inst_cellmath__45_0_I1630 (.Y(N5408), .A(inst_cellmath__25[42]), .B(inst_cellmath__25[41]));
NOR2XL inst_cellmath__45_0_I1631 (.Y(N5384), .A(N5408), .B(N5422));
NAND2XL inst_cellmath__45_0_I1632 (.Y(N5371), .A(inst_cellmath__25[44]), .B(inst_cellmath__25[43]));
NAND2XL inst_cellmath__45_0_I1633 (.Y(N5370), .A(inst_cellmath__25[46]), .B(inst_cellmath__25[45]));
NOR2XL inst_cellmath__45_0_I1634 (.Y(N5337), .A(N5371), .B(N5370));
NAND2BXL inst_cellmath__45_0_I1638 (.Y(N5338), .AN(inst_cellmath__45[0]), .B(inst_cellmath__25[25]));
NAND2BXL inst_cellmath__45_0_I1639 (.Y(N5361), .AN(N5373), .B(inst_cellmath__25[31]));
OR2XL inst_cellmath__45_0_I1640 (.Y(N5385), .A(N5403), .B(N5373));
NAND2BXL inst_cellmath__45_0_I1641 (.Y(N5333), .AN(N5373), .B(N5365));
NAND3BXL inst_cellmath__45_0_I1642 (.Y(N5351), .AN(N5373), .B(inst_cellmath__25[35]), .C(N5365));
OR2XL inst_cellmath__45_0_I1643 (.Y(N5394), .A(N5419), .B(N5373));
NAND2XL inst_cellmath__45_0_I1644 (.Y(N5344), .A(inst_cellmath__25[39]), .B(N5392));
NAND2BXL inst_cellmath__45_0_I1645 (.Y(N5404), .AN(N5422), .B(N5392));
NAND3BXL inst_cellmath__45_0_I1646 (.Y(N5369), .AN(N5422), .B(inst_cellmath__25[41]), .C(N5392));
NAND2XL inst_cellmath__45_0_I1647 (.Y(N5341), .A(N5384), .B(N5392));
NAND3XL inst_cellmath__45_0_I1648 (.Y(N5400), .A(inst_cellmath__25[43]), .B(N5384), .C(N5392));
NAND3BXL inst_cellmath__45_0_I1649 (.Y(N5366), .AN(N5371), .B(N5384), .C(N5392));
NAND4BXL inst_cellmath__45_0_I1650 (.Y(N5336), .AN(N5371), .B(inst_cellmath__25[45]), .C(N5392), .D(N5384));
NAND3XL hyperpropagate_4_1_A_I3712 (.Y(N8411), .A(N5337), .B(N5392), .C(N5384));
NOR2XL hyperpropagate_4_1_A_I3713 (.Y(inst_cellmath__45[24]), .A(inst_cellmath__25[47]), .B(N8411));
XNOR2X1 inst_cellmath__45_0_I1653 (.Y(inst_cellmath__45[1]), .A(inst_cellmath__45[0]), .B(inst_cellmath__25[25]));
XNOR2X1 inst_cellmath__45_0_I1654 (.Y(inst_cellmath__45[2]), .A(N5338), .B(inst_cellmath__25[26]));
XOR2XL inst_cellmath__45_0_I1655 (.Y(inst_cellmath__45[3]), .A(N5387), .B(inst_cellmath__25[27]));
XNOR2X1 inst_cellmath__45_0_I1656 (.Y(inst_cellmath__45[4]), .A(N5375), .B(inst_cellmath__25[28]));
XNOR2X1 inst_cellmath__45_0_I1657 (.Y(inst_cellmath__45[5]), .A(N5346), .B(inst_cellmath__25[29]));
XNOR2X1 inst_cellmath__45_0_I1658 (.Y(inst_cellmath__45[6]), .A(N5406), .B(inst_cellmath__25[30]));
XNOR2X1 inst_cellmath__45_0_I1659 (.Y(inst_cellmath__45[7]), .A(N5373), .B(inst_cellmath__25[31]));
XNOR2X1 inst_cellmath__45_0_I1660 (.Y(inst_cellmath__45[8]), .A(N5361), .B(inst_cellmath__25[32]));
XNOR2X1 inst_cellmath__45_0_I1661 (.Y(inst_cellmath__45[9]), .A(N5385), .B(inst_cellmath__25[33]));
XOR2XL inst_cellmath__45_0_I1662 (.Y(inst_cellmath__45[10]), .A(N5363), .B(inst_cellmath__25[34]));
XNOR2X1 inst_cellmath__45_0_I1663 (.Y(inst_cellmath__45[11]), .A(N5333), .B(inst_cellmath__25[35]));
XNOR2X1 inst_cellmath__45_0_I1664 (.Y(inst_cellmath__45[12]), .A(N5351), .B(inst_cellmath__25[36]));
XOR2XL inst_cellmath__45_0_I1665 (.Y(inst_cellmath__45[13]), .A(N5359), .B(inst_cellmath__25[37]));
XNOR2X1 inst_cellmath__45_0_I1666 (.Y(inst_cellmath__45[14]), .A(N5394), .B(inst_cellmath__25[38]));
XOR2XL inst_cellmath__45_0_I1667 (.Y(inst_cellmath__45[15]), .A(N5392), .B(inst_cellmath__25[39]));
XNOR2X1 inst_cellmath__45_0_I1668 (.Y(inst_cellmath__45[16]), .A(N5344), .B(inst_cellmath__25[40]));
XNOR2X1 inst_cellmath__45_0_I1669 (.Y(inst_cellmath__45[17]), .A(N5404), .B(inst_cellmath__25[41]));
XNOR2X1 inst_cellmath__45_0_I1670 (.Y(inst_cellmath__45[18]), .A(N5369), .B(inst_cellmath__25[42]));
XNOR2X1 inst_cellmath__45_0_I1671 (.Y(inst_cellmath__45[19]), .A(N5341), .B(inst_cellmath__25[43]));
XNOR2X1 inst_cellmath__45_0_I1672 (.Y(inst_cellmath__45[20]), .A(N5400), .B(inst_cellmath__25[44]));
XNOR2X1 inst_cellmath__45_0_I1673 (.Y(inst_cellmath__45[21]), .A(N5366), .B(inst_cellmath__25[45]));
XNOR2X1 inst_cellmath__45_0_I1674 (.Y(inst_cellmath__45[22]), .A(N5336), .B(inst_cellmath__25[46]));
NOR3BXL cynw_cm_float_mul_ieee_I1676 (.Y(inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
INVXL inst_cellmath__44__31__I1677 (.Y(N5500), .A(inst_cellmath__23));
AND2XL inst_cellmath__44__31__I1678 (.Y(N446), .A(inst_cellmath__5), .B(N5500));
NOR3BXL cynw_cm_float_mul_ieee_I1679 (.Y(inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
AND2XL cynw_cm_float_mul_ieee_I1680 (.Y(N445), .A(inst_cellmath__6), .B(inst_cellmath__23));
NOR3BXL cynw_cm_float_mul_ieee_I1681 (.Y(inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3XL cynw_cm_float_mul_ieee_I1682 (.Y(inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
NOR2XL inst_cellmath__34_0_I1683 (.Y(N5536), .A(inst_cellmath__25[19]), .B(inst_cellmath__25[17]));
NOR2XL inst_cellmath__34_0_I1684 (.Y(N5547), .A(inst_cellmath__25[15]), .B(inst_cellmath__25[13]));
NOR2XL inst_cellmath__34_0_I1687 (.Y(N5530), .A(inst_cellmath__25[3]), .B(inst_cellmath__25[22]));
NOR2XL inst_cellmath__34_0_I1688 (.Y(N5540), .A(inst_cellmath__25[20]), .B(inst_cellmath__25[18]));
NAND2XL inst_cellmath__34_0_I1693 (.Y(N5545), .A(N5536), .B(N5547));
OR4X1 inst_cellmath__34_0_I10208 (.Y(N5554), .A(inst_cellmath__25[5]), .B(inst_cellmath__25[9]), .C(inst_cellmath__25[7]), .D(inst_cellmath__25[11]));
OR4X1 inst_cellmath__34_0_I10209 (.Y(N5528), .A(inst_cellmath__25[10]), .B(inst_cellmath__25[14]), .C(inst_cellmath__25[12]), .D(inst_cellmath__25[16]));
OR4X1 inst_cellmath__34_0_I10210 (.Y(N5538), .A(inst_cellmath__25[2]), .B(inst_cellmath__25[6]), .C(inst_cellmath__25[4]), .D(inst_cellmath__25[8]));
NOR4X1 inst_cellmath__34_0_I1697 (.Y(N5558), .A(inst_cellmath__25[0]), .B(inst_cellmath__25[1]), .C(inst_cellmath__25[21]), .D(N5545));
NOR2XL inst_cellmath__34_0_I1698 (.Y(N5552), .A(N5528), .B(N5538));
NAND3XL inst_cellmath__34_0_I1699 (.Y(N5532), .A(N5530), .B(N5540), .C(N5558));
NOR2XL inst_cellmath__34_0_I1700 (.Y(N5543), .A(N5554), .B(N5532));
NAND2XL inst_cellmath__34_0_I1701 (.Y(inst_cellmath__34), .A(N5552), .B(N5543));
OA21X1 cynw_cm_float_mul_ieee_I3663 (.Y(N444), .A0(inst_cellmath__25[24]), .A1(inst_cellmath__34), .B0(inst_cellmath__4));
OR4X1 cynw_cm_float_mul_ieee_I1704 (.Y(N447), .A(inst_cellmath__8), .B(N445), .C(N446), .D(N444));
OAI21XL cynw_cm_float_mul_ieee_I3664 (.Y(N450), .A0(N445), .A1(N446), .B0(inst_cellmath__34));
OAI2BB1X1 cynw_cm_float_mul_ieee_I3665 (.Y(inst_cellmath__44), .A0N(inst_cellmath__25[23]), .A1N(N447), .B0(N450));
AOI21X1 cynw_cm_float_mul_ieee_I3667 (.Y(inst_cellmath__38), .A0(inst_cellmath__45[24]), .A1(inst_cellmath__44), .B0(inst_cellmath__24[47]));
INVXL inst_cellmath__30_0_I1711 (.Y(N5627), .A(a_exp[7]));
XNOR2X1 inst_cellmath__30_0_I1712 (.Y(inst_cellmath__30[0]), .A(b_exp[0]), .B(a_exp[0]));
OR2XL inst_cellmath__30_0_I1713 (.Y(N5631), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 inst_cellmath__30_0_I1714 (.CO(N5624), .S(inst_cellmath__30[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(N5631));
ADDFX1 inst_cellmath__30_0_I1715 (.CO(N5643), .S(inst_cellmath__30[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(N5624));
ADDFX1 inst_cellmath__30_0_I1716 (.CO(N5655), .S(inst_cellmath__30[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(N5643));
ADDFX1 inst_cellmath__30_0_I1717 (.CO(N5637), .S(inst_cellmath__30[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(N5655));
ADDFX1 inst_cellmath__30_0_I1718 (.CO(N5652), .S(inst_cellmath__30[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(N5637));
ADDFX1 inst_cellmath__30_0_I1719 (.CO(N5632), .S(inst_cellmath__30[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(N5652));
ADDFX1 inst_cellmath__30_0_I1720 (.CO(N5647), .S(inst_cellmath__30[7]), .A(N5627), .B(b_exp[7]), .CI(N5632));
XNOR2X1 inst_cellmath__30_0_I1721 (.Y(inst_cellmath__30[8]), .A(a_exp[7]), .B(N5647));
NOR2XL inst_cellmath__30_0_I1722 (.Y(inst_cellmath__30[9]), .A(a_exp[7]), .B(N5647));
INVXL inst_cellmath__31_0_I1723 (.Y(inst_cellmath__31[0]), .A(inst_cellmath__30[0]));
NOR2BX1 inst_cellmath__31_0_I1724 (.Y(N5697), .AN(inst_cellmath__30[1]), .B(inst_cellmath__31[0]));
AND2XL inst_cellmath__31_0_I1725 (.Y(N5682), .A(inst_cellmath__30[2]), .B(N5697));
XNOR2X1 inst_cellmath__31_0_I1726 (.Y(inst_cellmath__31[1]), .A(inst_cellmath__31[0]), .B(inst_cellmath__30[1]));
XOR2XL inst_cellmath__31_0_I1727 (.Y(inst_cellmath__31[2]), .A(N5697), .B(inst_cellmath__30[2]));
AND2XL inst_cellmath__31_0_I1728 (.Y(N5701), .A(inst_cellmath__30[3]), .B(N5682));
AND3XL inst_cellmath__31_0_I1729 (.Y(N5700), .A(inst_cellmath__30[4]), .B(inst_cellmath__30[5]), .C(N5701));
AND3XL inst_cellmath__31_0_I1730 (.Y(N5691), .A(inst_cellmath__30[6]), .B(inst_cellmath__30[7]), .C(N5700));
NAND2XL inst_cellmath__31_0_I1731 (.Y(N5681), .A(inst_cellmath__30[4]), .B(N5701));
NAND2XL inst_cellmath__31_0_I1732 (.Y(N5699), .A(inst_cellmath__30[6]), .B(N5700));
NAND2XL inst_cellmath__31_0_I1733 (.Y(N5690), .A(inst_cellmath__30[8]), .B(N5691));
XOR2XL inst_cellmath__31_0_I1734 (.Y(inst_cellmath__31[3]), .A(N5682), .B(inst_cellmath__30[3]));
XOR2XL inst_cellmath__31_0_I1735 (.Y(inst_cellmath__31[4]), .A(N5701), .B(inst_cellmath__30[4]));
XNOR2X1 inst_cellmath__31_0_I1736 (.Y(inst_cellmath__31[5]), .A(N5681), .B(inst_cellmath__30[5]));
XOR2XL inst_cellmath__31_0_I1737 (.Y(inst_cellmath__31[6]), .A(N5700), .B(inst_cellmath__30[6]));
XNOR2X1 inst_cellmath__31_0_I1738 (.Y(inst_cellmath__31[7]), .A(N5699), .B(inst_cellmath__30[7]));
XOR2XL inst_cellmath__31_0_I1739 (.Y(inst_cellmath__31[8]), .A(N5691), .B(inst_cellmath__30[8]));
XNOR2X1 inst_cellmath__31_0_I1740 (.Y(inst_cellmath__31[9]), .A(N5690), .B(inst_cellmath__30[9]));
MX2XL inst_cellmath__48_0_I1741 (.Y(inst_cellmath__48[0]), .A(inst_cellmath__31[0]), .B(inst_cellmath__30[0]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1742 (.Y(inst_cellmath__48[1]), .A(inst_cellmath__31[1]), .B(inst_cellmath__30[1]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1743 (.Y(inst_cellmath__48[2]), .A(inst_cellmath__31[2]), .B(inst_cellmath__30[2]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1744 (.Y(inst_cellmath__48[3]), .A(inst_cellmath__31[3]), .B(inst_cellmath__30[3]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1745 (.Y(inst_cellmath__48[4]), .A(inst_cellmath__31[4]), .B(inst_cellmath__30[4]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1746 (.Y(inst_cellmath__48[5]), .A(inst_cellmath__31[5]), .B(inst_cellmath__30[5]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1747 (.Y(inst_cellmath__48[6]), .A(inst_cellmath__31[6]), .B(inst_cellmath__30[6]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1748 (.Y(inst_cellmath__48[7]), .A(inst_cellmath__31[7]), .B(inst_cellmath__30[7]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1749 (.Y(inst_cellmath__48[8]), .A(inst_cellmath__31[8]), .B(inst_cellmath__30[8]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1750 (.Y(inst_cellmath__48[9]), .A(inst_cellmath__31[9]), .B(inst_cellmath__30[9]), .S0(inst_cellmath__38));
NAND2XL inst_cellmath__51__49__I1751 (.Y(N5768), .A(inst_cellmath__48[1]), .B(inst_cellmath__48[6]));
NAND2XL inst_cellmath__51__49__I1752 (.Y(N5772), .A(inst_cellmath__48[0]), .B(inst_cellmath__48[5]));
NAND2XL inst_cellmath__51__49__I1753 (.Y(N5775), .A(inst_cellmath__48[4]), .B(inst_cellmath__48[2]));
NAND2XL inst_cellmath__51__49__I1754 (.Y(N5763), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[3]));
NOR4X1 inst_cellmath__51__49__I3688 (.Y(N461), .A(N5768), .B(N5763), .C(N5775), .D(N5772));
NOR2XL andori2bb1_A_I3714 (.Y(N8417), .A(inst_cellmath__48[8]), .B(N461));
NOR2XL andori2bb1_A_I3715 (.Y(inst_cellmath__51), .A(N8417), .B(inst_cellmath__48[9]));
NAND2XL cynw_cm_float_mul_ieee_I1760 (.Y(inst_cellmath__28), .A(inst_cellmath__20), .B(inst_cellmath__13));
NAND2XL cynw_cm_float_mul_ieee_I1761 (.Y(inst_cellmath__27), .A(inst_cellmath__21), .B(inst_cellmath__14));
NOR2XL inst_cellmath__50__50__I1762 (.Y(N5813), .A(inst_cellmath__48[8]), .B(inst_cellmath__48[1]));
NOR2XL inst_cellmath__50__50__I1763 (.Y(N5801), .A(inst_cellmath__48[6]), .B(inst_cellmath__48[9]));
NAND2XL inst_cellmath__50__50__I1764 (.Y(N5815), .A(N5813), .B(N5801));
NOR4X1 inst_cellmath__50__50__I1765 (.Y(N5812), .A(inst_cellmath__48[0]), .B(inst_cellmath__48[2]), .C(inst_cellmath__48[4]), .D(inst_cellmath__48[5]));
NOR3XL inst_cellmath__50__50__I1766 (.Y(N5808), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[3]), .C(N5815));
NOR4X1 inst_cellmath__49_1_I1768 (.Y(N5830), .A(inst_cellmath__28), .B(inst_cellmath__27), .C(inst_cellmath__26), .D(inst_cellmath__48[9]));
OAI2BB1X1 inst_cellmath__49_1_I3671 (.Y(N5823), .A0N(N5812), .A1N(N5808), .B0(N5830));
OR2XL inst_cellmath__49_1_I1770 (.Y(inst_cellmath__49), .A(N5823), .B(inst_cellmath__51));
OR2XL cynw_cm_float_mul_ieee_I1771 (.Y(N470), .A(inst_cellmath__27), .B(inst_cellmath__26));
OR2XL cynw_cm_float_mul_ieee_I1772 (.Y(N442), .A(inst_cellmath__30[8]), .B(inst_cellmath__30[7]));
NAND2BXL cynw_cm_float_mul_ieee_I1773 (.Y(inst_cellmath__32), .AN(inst_cellmath__30[9]), .B(N442));
NOR2XL cynw_cm_float_mul_ieee_I1774 (.Y(N469), .A(inst_cellmath__28), .B(inst_cellmath__32));
NAND2XL inst_cellmath__7_0_I1775 (.Y(N5852), .A(rm[0]), .B(rm[1]));
NOR2XL inst_cellmath__7_0_I1776 (.Y(inst_cellmath__7), .A(rm[2]), .B(N5852));
MXI2XL inst_cellmath__42_0_I1778 (.Y(N5860), .A(inst_cellmath__7), .B(N5500), .S0(inst_cellmath__6));
MX2XL inst_cellmath__42_0_I1779 (.Y(inst_cellmath__42), .A(N5860), .B(N5500), .S0(inst_cellmath__5));
AOI21XL inst_cellmath__52_0_I1781 (.Y(N5893), .A0(inst_cellmath__42), .A1(N469), .B0(N470));
OR2XL inst_cellmath__52_0_I1782 (.Y(N5874), .A(N469), .B(N470));
INVXL inst_cellmath__52_0_I1783 (.Y(N5870), .A(inst_cellmath__48[0]));
INVXL inst_cellmath__52_0_I1784 (.Y(N5887), .A(inst_cellmath__49));
INVXL inst_cellmath__52_0_I1785 (.Y(N5884), .A(N5887));
MXI2XL inst_cellmath__52_0_I1786 (.Y(x[23]), .A(N5870), .B(N5893), .S0(N5884));
MX2XL inst_cellmath__52_0_I1787 (.Y(x[24]), .A(inst_cellmath__48[1]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1788 (.Y(x[25]), .A(inst_cellmath__48[2]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1789 (.Y(x[26]), .A(inst_cellmath__48[3]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1790 (.Y(x[27]), .A(inst_cellmath__48[4]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1791 (.Y(x[28]), .A(inst_cellmath__48[5]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1792 (.Y(x[29]), .A(inst_cellmath__48[6]), .B(N5874), .S0(N5884));
MX2XL inst_cellmath__52_0_I1793 (.Y(x[30]), .A(inst_cellmath__48[7]), .B(N5874), .S0(N5884));
OR4X1 inst_cellmath__47_0_I1794 (.Y(N5914), .A(inst_cellmath__28), .B(inst_cellmath__27), .C(inst_cellmath__26), .D(inst_cellmath__42));
NOR2XL inst_cellmath__47_0_I1795 (.Y(inst_cellmath__47), .A(N5914), .B(inst_cellmath__32));
NOR2XL inst_cellmath__53_U_I1796 (.Y(N5925), .A(inst_cellmath__26), .B(inst_cellmath__47));
MXI2XL inst_cellmath__53_U_I1797 (.Y(N5923), .A(inst_cellmath__25[46]), .B(inst_cellmath__45[22]), .S0(inst_cellmath__44));
MXI2XL inst_cellmath__53_U_I1798 (.Y(x[22]), .A(N5923), .B(N5925), .S0(inst_cellmath__49));
NOR2X1 inst_cellmath__53_M_I3673 (.Y(N8378), .A(inst_cellmath__26), .B(N5887));
NAND3BXL inst_cellmath__53_M_I1801 (.Y(N6014), .AN(inst_cellmath__15), .B(inst_cellmath__22), .C(inst_cellmath__26));
NOR2X1 inst_cellmath__53_M_I3675 (.Y(N8380), .A(N6014), .B(N5887));
NAND2XL inst_cellmath__53_M_I1803 (.Y(N6095), .A(inst_cellmath__15), .B(inst_cellmath__26));
NOR2X1 inst_cellmath__53_M_I3677 (.Y(N8382), .A(N6095), .B(N5887));
NOR2BX1 inst_cellmath__53_M_I1805 (.Y(N5987), .AN(N5887), .B(inst_cellmath__44));
AND2XL inst_cellmath__53_M_I1806 (.Y(N6028), .A(inst_cellmath__44), .B(N5887));
AOI22XL inst_cellmath__53_M_I1807 (.Y(N6114), .A0(inst_cellmath__45[0]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[24]));
AOI22XL inst_cellmath__53_M_I1808 (.Y(N6008), .A0(inst_cellmath__45[1]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[25]));
AOI22XL inst_cellmath__53_M_I1809 (.Y(N6088), .A0(inst_cellmath__45[2]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[26]));
AOI22XL inst_cellmath__53_M_I1810 (.Y(N5982), .A0(inst_cellmath__45[3]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[27]));
AOI22XL inst_cellmath__53_M_I1811 (.Y(N6066), .A0(inst_cellmath__45[4]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[28]));
AOI22XL inst_cellmath__53_M_I1812 (.Y(N5957), .A0(inst_cellmath__45[5]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[29]));
AOI22XL inst_cellmath__53_M_I1813 (.Y(N6040), .A0(inst_cellmath__45[6]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[30]));
AOI22XL inst_cellmath__53_M_I1814 (.Y(N5933), .A0(inst_cellmath__45[7]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[31]));
AOI22XL inst_cellmath__53_M_I1815 (.Y(N6018), .A0(inst_cellmath__45[8]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[32]));
AOI22XL inst_cellmath__53_M_I1816 (.Y(N6100), .A0(inst_cellmath__45[9]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[33]));
AOI22XL inst_cellmath__53_M_I1817 (.Y(N5992), .A0(inst_cellmath__45[10]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[34]));
AOI22XL inst_cellmath__53_M_I1818 (.Y(N6077), .A0(inst_cellmath__45[11]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[35]));
AOI22XL inst_cellmath__53_M_I1819 (.Y(N5967), .A0(inst_cellmath__45[12]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[36]));
AOI22XL inst_cellmath__53_M_I1820 (.Y(N6051), .A0(inst_cellmath__45[13]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[37]));
AOI22XL inst_cellmath__53_M_I1821 (.Y(N5941), .A0(inst_cellmath__45[14]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[38]));
AOI22XL inst_cellmath__53_M_I1822 (.Y(N6027), .A0(inst_cellmath__45[15]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[39]));
AOI22XL inst_cellmath__53_M_I1823 (.Y(N6109), .A0(inst_cellmath__45[16]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[40]));
AOI22XL inst_cellmath__53_M_I1824 (.Y(N6002), .A0(inst_cellmath__45[17]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[41]));
AOI22XL inst_cellmath__53_M_I1825 (.Y(N6084), .A0(inst_cellmath__45[18]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[42]));
AOI22XL inst_cellmath__53_M_I1826 (.Y(N5977), .A0(inst_cellmath__45[19]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[43]));
AOI22XL inst_cellmath__53_M_I1827 (.Y(N6061), .A0(inst_cellmath__45[20]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[44]));
AOI22XL inst_cellmath__53_M_I1828 (.Y(N5951), .A0(inst_cellmath__45[21]), .A1(N6028), .B0(N5987), .B1(inst_cellmath__25[45]));
AOI22XL inst_cellmath__53_M_I1829 (.Y(N5984), .A0(b_man[0]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1830 (.Y(N5959), .A0(b_man[1]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1831 (.Y(N5934), .A0(b_man[2]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1832 (.Y(N6102), .A0(b_man[3]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1833 (.Y(N6079), .A0(b_man[4]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1834 (.Y(N6053), .A0(b_man[5]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1835 (.Y(N6030), .A0(b_man[6]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1836 (.Y(N6004), .A0(b_man[7]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1837 (.Y(N5978), .A0(b_man[8]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1838 (.Y(N5953), .A0(b_man[9]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1839 (.Y(N5930), .A0(b_man[10]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1840 (.Y(N6096), .A0(b_man[11]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1841 (.Y(N6073), .A0(b_man[12]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1842 (.Y(N6047), .A0(b_man[13]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1843 (.Y(N6024), .A0(b_man[14]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1844 (.Y(N5999), .A0(b_man[15]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1845 (.Y(N5973), .A0(b_man[16]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1846 (.Y(N5948), .A0(b_man[17]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1847 (.Y(N6117), .A0(b_man[18]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1848 (.Y(N6091), .A0(b_man[19]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1849 (.Y(N6069), .A0(b_man[20]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1850 (.Y(N6043), .A0(b_man[21]), .A1(N8380), .B0(N8378), .B1(inst_cellmath__47));
NAND2XL inst_cellmath__53_M_I1851 (.Y(N6020), .A(N8382), .B(a_man[0]));
NAND2XL inst_cellmath__53_M_I1852 (.Y(N6104), .A(N8382), .B(a_man[1]));
NAND2XL inst_cellmath__53_M_I1853 (.Y(N5996), .A(N8382), .B(a_man[2]));
NAND2XL inst_cellmath__53_M_I1854 (.Y(N6080), .A(N8382), .B(a_man[3]));
NAND2XL inst_cellmath__53_M_I1855 (.Y(N5970), .A(N8382), .B(a_man[4]));
NAND2XL inst_cellmath__53_M_I1856 (.Y(N6055), .A(N8382), .B(a_man[5]));
NAND2XL inst_cellmath__53_M_I1857 (.Y(N5943), .A(N8382), .B(a_man[6]));
NAND2XL inst_cellmath__53_M_I1858 (.Y(N6032), .A(N8382), .B(a_man[7]));
NAND2XL inst_cellmath__53_M_I1859 (.Y(N6112), .A(N8382), .B(a_man[8]));
NAND2XL inst_cellmath__53_M_I1860 (.Y(N6005), .A(N8382), .B(a_man[9]));
NAND2XL inst_cellmath__53_M_I1861 (.Y(N6086), .A(N8382), .B(a_man[10]));
NAND2XL inst_cellmath__53_M_I1862 (.Y(N5980), .A(N8382), .B(a_man[11]));
NAND2XL inst_cellmath__53_M_I1863 (.Y(N6063), .A(N8382), .B(a_man[12]));
NAND2XL inst_cellmath__53_M_I1864 (.Y(N5955), .A(N8382), .B(a_man[13]));
NAND2XL inst_cellmath__53_M_I1865 (.Y(N6038), .A(N8382), .B(a_man[14]));
NAND2XL inst_cellmath__53_M_I1866 (.Y(N5931), .A(N8382), .B(a_man[15]));
NAND2XL inst_cellmath__53_M_I1867 (.Y(N6016), .A(N8382), .B(a_man[16]));
NAND2XL inst_cellmath__53_M_I1868 (.Y(N6098), .A(N8382), .B(a_man[17]));
NAND2XL inst_cellmath__53_M_I1869 (.Y(N5990), .A(N8382), .B(a_man[18]));
NAND2XL inst_cellmath__53_M_I1870 (.Y(N6075), .A(N8382), .B(a_man[19]));
NAND2XL inst_cellmath__53_M_I1871 (.Y(N5965), .A(N8382), .B(a_man[20]));
NAND2XL inst_cellmath__53_M_I1872 (.Y(N6048), .A(N8382), .B(a_man[21]));
NAND3XL inst_cellmath__53_M_I1873 (.Y(x[0]), .A(N6020), .B(N6114), .C(N5984));
NAND3XL inst_cellmath__53_M_I1874 (.Y(x[1]), .A(N6104), .B(N6008), .C(N5959));
NAND3XL inst_cellmath__53_M_I1875 (.Y(x[2]), .A(N5996), .B(N6088), .C(N5934));
NAND3XL inst_cellmath__53_M_I1876 (.Y(x[3]), .A(N6080), .B(N5982), .C(N6102));
NAND3XL inst_cellmath__53_M_I1877 (.Y(x[4]), .A(N5970), .B(N6066), .C(N6079));
NAND3XL inst_cellmath__53_M_I1878 (.Y(x[5]), .A(N6055), .B(N5957), .C(N6053));
NAND3XL inst_cellmath__53_M_I1879 (.Y(x[6]), .A(N5943), .B(N6040), .C(N6030));
NAND3XL inst_cellmath__53_M_I1880 (.Y(x[7]), .A(N6032), .B(N5933), .C(N6004));
NAND3XL inst_cellmath__53_M_I1881 (.Y(x[8]), .A(N6112), .B(N6018), .C(N5978));
NAND3XL inst_cellmath__53_M_I1882 (.Y(x[9]), .A(N6005), .B(N6100), .C(N5953));
NAND3XL inst_cellmath__53_M_I1883 (.Y(x[10]), .A(N6086), .B(N5992), .C(N5930));
NAND3XL inst_cellmath__53_M_I1884 (.Y(x[11]), .A(N5980), .B(N6077), .C(N6096));
NAND3XL inst_cellmath__53_M_I1885 (.Y(x[12]), .A(N6063), .B(N5967), .C(N6073));
NAND3XL inst_cellmath__53_M_I1886 (.Y(x[13]), .A(N5955), .B(N6051), .C(N6047));
NAND3XL inst_cellmath__53_M_I1887 (.Y(x[14]), .A(N6038), .B(N5941), .C(N6024));
NAND3XL inst_cellmath__53_M_I1888 (.Y(x[15]), .A(N5931), .B(N6027), .C(N5999));
NAND3XL inst_cellmath__53_M_I1889 (.Y(x[16]), .A(N6016), .B(N6109), .C(N5973));
NAND3XL inst_cellmath__53_M_I1890 (.Y(x[17]), .A(N6098), .B(N6002), .C(N5948));
NAND3XL inst_cellmath__53_M_I1891 (.Y(x[18]), .A(N5990), .B(N6084), .C(N6117));
NAND3XL inst_cellmath__53_M_I1892 (.Y(x[19]), .A(N6075), .B(N5977), .C(N6091));
NAND3XL inst_cellmath__53_M_I1893 (.Y(x[20]), .A(N5965), .B(N6061), .C(N6069));
NAND3XL inst_cellmath__53_M_I1894 (.Y(x[21]), .A(N6048), .B(N5951), .C(N6043));
assign inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  urfzSw/Wqh8= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



