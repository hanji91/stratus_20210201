/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:07:19 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_3 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
wire  inst_cellmath__5,
	inst_cellmath__6,
	inst_cellmath__7,
	inst_cellmath__8,
	inst_cellmath__10,
	inst_cellmath__12,
	inst_cellmath__13,
	inst_cellmath__14,
	inst_cellmath__15,
	inst_cellmath__17,
	inst_cellmath__19,
	inst_cellmath__20,
	inst_cellmath__21,
	inst_cellmath__22,
	inst_cellmath__23;
wire [47:0] inst_cellmath__24,
	inst_cellmath__25;
wire  inst_cellmath__26,
	inst_cellmath__27,
	inst_cellmath__28;
wire [9:0] inst_cellmath__30,
	inst_cellmath__31;
wire  inst_cellmath__32,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42,
	inst_cellmath__44;
wire [24:0] inst_cellmath__45;
wire  inst_cellmath__47;
wire [9:0] inst_cellmath__48;
wire  inst_cellmath__49,
	inst_cellmath__51;
wire N440,N441,N442,N443,N444,N445,N446 
	,N447,N450,N461,N469,N470,N1896,N1898,N1919 
	,N1927,N1930,N1932,N1936,N1938,N1941,N1947,N1951 
	,N1976,N1981,N1985,N1988,N2007,N2009,N2030,N2038 
	,N2041,N2043,N2047,N2049,N2052,N2058,N2062,N2087 
	,N2092,N2096,N2099,N2131,N2136,N2143,N2144,N2145 
	,N2146,N2147,N2148,N2149,N2150,N2151,N2152,N2153 
	,N2154,N2155,N2156,N2157,N2158,N2159,N2160,N2161 
	,N2162,N2163,N2164,N2165,N2166,N2168,N2169,N2170 
	,N2171,N2172,N2173,N2174,N2175,N2176,N2177,N2179 
	,N2180,N2181,N2182,N2183,N2185,N2186,N2187,N2188 
	,N2189,N2190,N2191,N2192,N2193,N2194,N2195,N2196 
	,N2197,N2198,N2199,N2200,N2201,N2202,N2203,N2204 
	,N2205,N2206,N2207,N2208,N2209,N2210,N2211,N2212 
	,N2213,N2214,N2215,N2216,N2217,N2218,N2219,N2220 
	,N2221,N2222,N2223,N2224,N2225,N2227,N2228,N2230 
	,N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238 
	,N2239,N2240,N2241,N2244,N2245,N2246,N2247,N2248 
	,N2249,N2250,N2252,N2253,N2254,N2255,N2256,N2257 
	,N2258,N2259,N2260,N2261,N2262,N2263,N2264,N2265 
	,N2266,N2267,N2268,N2269,N2270,N2271,N2272,N2273 
	,N2274,N2275,N2276,N2277,N2278,N2279,N2280,N2282 
	,N2283,N2284,N2285,N2286,N2287,N2288,N2289,N2290 
	,N2291,N2292,N2293,N2294,N2295,N2296,N2297,N2298 
	,N2299,N2300,N2301,N2302,N2304,N2306,N2307,N2308 
	,N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316 
	,N2317,N2318,N2319,N2320,N2321,N2322,N2324,N2325 
	,N2326,N2327,N2328,N2329,N2330,N2331,N2332,N2333 
	,N2334,N2335,N2336,N2337,N2338,N2340,N2341,N2342 
	,N2343,N2344,N2345,N2346,N2347,N2348,N2349,N2350 
	,N2351,N2352,N2353,N2354,N2355,N2356,N2357,N2358 
	,N2359,N2360,N2361,N2362,N2363,N2364,N2366,N2367 
	,N2368,N2369,N2370,N2372,N2373,N2374,N2375,N2376 
	,N2377,N2378,N2379,N2380,N2381,N2382,N2383,N2384 
	,N2385,N2387,N2388,N2389,N2390,N2391,N2392,N2393 
	,N2394,N2396,N2397,N2398,N2399,N2400,N2401,N2402 
	,N2403,N2404,N2405,N2406,N2407,N2408,N2409,N2410 
	,N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2418 
	,N2419,N2420,N2421,N2422,N2423,N2424,N2425,N2426 
	,N2427,N2428,N2429,N2431,N2432,N2433,N2435,N2436 
	,N2437,N2438,N2439,N2440,N2441,N2442,N2443,N2444 
	,N2446,N2447,N2448,N2449,N2450,N2451,N2452,N2453 
	,N2454,N2455,N2456,N2457,N2459,N2460,N2461,N2462 
	,N2463,N2464,N2465,N2466,N2467,N2468,N2469,N2470 
	,N2471,N2472,N2473,N2474,N2476,N2477,N2478,N2479 
	,N2480,N2481,N2482,N2483,N2484,N2485,N2486,N2487 
	,N2488,N2489,N2491,N2492,N2493,N2494,N2495,N2496 
	,N2497,N2498,N2499,N2500,N2501,N2502,N2503,N2504 
	,N2505,N2506,N2507,N2508,N2509,N2510,N2511,N2512 
	,N2514,N2515,N2516,N2517,N2518,N2520,N2521,N2522 
	,N2524,N2525,N2526,N2527,N2528,N2529,N2530,N2531 
	,N2532,N2533,N2534,N2535,N2536,N2537,N2539,N2540 
	,N2541,N2542,N2543,N2544,N2545,N2546,N2547,N2548 
	,N2549,N2550,N2551,N2552,N2553,N2554,N2555,N2556 
	,N2557,N2558,N2559,N2560,N2561,N2562,N2563,N2564 
	,N2565,N2566,N2567,N2568,N2569,N2570,N2571,N2572 
	,N2573,N2574,N2575,N2576,N2577,N2579,N2580,N2582 
	,N2583,N2584,N2585,N2586,N2587,N2588,N2589,N2590 
	,N2591,N2592,N2593,N2594,N2595,N2596,N2597,N2598 
	,N2600,N2601,N2602,N2603,N2604,N2606,N2607,N2608 
	,N2609,N2610,N2611,N2612,N2613,N2614,N2615,N2616 
	,N2617,N2618,N2619,N2620,N2621,N2622,N2623,N2624 
	,N2625,N2626,N2627,N2628,N2629,N2630,N2631,N2632 
	,N2633,N2634,N2635,N2636,N2638,N2639,N2640,N2641 
	,N2642,N2644,N2645,N2646,N2647,N2649,N2650,N2651 
	,N2652,N2653,N2654,N2655,N2656,N2657,N2658,N2659 
	,N2660,N2661,N2662,N2663,N2664,N2666,N2667,N2668 
	,N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676 
	,N2677,N2678,N2679,N2680,N2681,N2682,N2683,N2685 
	,N2686,N2687,N2688,N2689,N2690,N2691,N2692,N2693 
	,N2694,N2695,N2696,N2697,N2698,N2700,N2701,N2702 
	,N2703,N2704,N2705,N2706,N2707,N2708,N2709,N2710 
	,N2711,N2712,N2713,N2714,N2715,N2716,N2717,N2718 
	,N2719,N2720,N2721,N2722,N2723,N2724,N2725,N2726 
	,N2727,N2728,N2729,N2730,N2731,N2732,N2734,N2736 
	,N2737,N2738,N2739,N2740,N2741,N2742,N2743,N2744 
	,N2745,N2746,N2747,N2748,N2749,N2751,N2752,N2753 
	,N2754,N2755,N2756,N2757,N2758,N2759,N2760,N2761 
	,N2762,N2763,N2764,N2765,N2766,N2767,N2768,N2769 
	,N2770,N2771,N2772,N2773,N2774,N2775,N2776,N2777 
	,N2778,N2779,N2780,N2781,N2782,N2783,N2784,N2785 
	,N2786,N2787,N2788,N2789,N2790,N2791,N2792,N2793 
	,N2794,N2796,N2797,N2798,N2799,N2800,N2801,N2802 
	,N2803,N2804,N2805,N2806,N2807,N2808,N2809,N2811 
	,N2812,N2813,N2814,N2816,N2817,N2818,N2819,N2820 
	,N2821,N2822,N2823,N2824,N2825,N2826,N2827,N2828 
	,N2829,N2830,N2831,N2832,N2833,N2834,N2835,N2836 
	,N2837,N2838,N2839,N2840,N2841,N2842,N2843,N2844 
	,N2845,N2846,N2847,N2848,N2849,N2851,N2852,N2853 
	,N2855,N2856,N2857,N2858,N2859,N2860,N2861,N2862 
	,N2863,N2864,N2865,N2866,N2867,N2868,N2869,N2870 
	,N2871,N2872,N2873,N2874,N2876,N2877,N2878,N2879 
	,N2880,N2881,N2882,N2883,N2884,N2885,N2886,N2887 
	,N2888,N2889,N2890,N2891,N2892,N2893,N2894,N2895 
	,N2897,N2898,N2899,N2900,N2901,N2902,N2903,N2904 
	,N2905,N2906,N2907,N2908,N2909,N2910,N2911,N2912 
	,N2913,N2914,N2915,N2916,N2917,N2918,N2919,N2920 
	,N2921,N2922,N2923,N2924,N2925,N2926,N2927,N2928 
	,N2929,N2930,N2931,N2932,N2933,N2934,N2935,N2936 
	,N2937,N2939,N2940,N2941,N2942,N2944,N2945,N2946 
	,N2947,N2948,N2949,N2950,N2951,N2952,N2953,N2954 
	,N2955,N2956,N2958,N2959,N2960,N2961,N2962,N2963 
	,N2964,N2965,N2966,N2968,N2969,N2970,N2971,N2972 
	,N2973,N2974,N2975,N2976,N2977,N2978,N2979,N2980 
	,N2981,N2982,N2983,N2984,N2985,N2986,N2987,N2988 
	,N2989,N2990,N2991,N2992,N2993,N2994,N2995,N2996 
	,N2997,N2998,N2999,N3000,N3001,N3002,N3003,N3005 
	,N3006,N3007,N3008,N3009,N3010,N3011,N3012,N3013 
	,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021 
	,N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029 
	,N3030,N3031,N3032,N3034,N3035,N3036,N3037,N3038 
	,N3039,N3040,N3041,N3042,N3043,N3044,N3045,N3046 
	,N3047,N3048,N3050,N3051,N3052,N3053,N3054,N3055 
	,N3056,N3057,N3058,N3059,N3060,N3061,N3063,N3064 
	,N3065,N3066,N3067,N3068,N3069,N3070,N3071,N3072 
	,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080 
	,N3081,N3082,N3083,N3084,N3085,N3086,N3087,N3088 
	,N3090,N3091,N3092,N3093,N3094,N3095,N3096,N3097 
	,N3098,N3099,N3100,N3101,N3102,N3103,N3104,N3105 
	,N3107,N3108,N3109,N3110,N3111,N3112,N3113,N3114 
	,N3115,N3116,N3117,N3118,N3119,N3120,N3121,N3122 
	,N3123,N3124,N3125,N3126,N3127,N3128,N3129,N3130 
	,N3131,N3132,N3133,N3134,N3135,N3136,N3137,N3138 
	,N3139,N3140,N3141,N3142,N3143,N3144,N3146,N3147 
	,N3148,N3149,N3150,N3152,N3153,N3154,N3155,N3156 
	,N3157,N3158,N3159,N3160,N3161,N3162,N3163,N3164 
	,N3166,N3167,N3168,N3169,N3170,N3171,N3172,N3174 
	,N3175,N3176,N3177,N3178,N3179,N3180,N3181,N3182 
	,N3183,N3184,N3185,N3186,N3187,N3188,N3189,N3190 
	,N3191,N3192,N3193,N3194,N3195,N3196,N3197,N3198 
	,N3199,N3200,N3201,N3202,N3203,N3204,N3206,N3207 
	,N3208,N3209,N3210,N3211,N3212,N3213,N3214,N3215 
	,N3216,N3217,N3218,N3219,N3220,N3221,N3222,N3223 
	,N3224,N3225,N3226,N3227,N3228,N3229,N3230,N3231 
	,N3233,N3234,N3235,N3236,N3237,N3238,N3239,N3240 
	,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3249 
	,N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257 
	,N3258,N3259,N3260,N3261,N3262,N3263,N3264,N3265 
	,N3266,N3267,N3268,N3269,N3270,N3271,N3272,N3273 
	,N3274,N3275,N3276,N3277,N3278,N3279,N3280,N3281 
	,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289 
	,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298 
	,N3299,N3300,N3301,N3302,N3303,N3304,N3305,N3306 
	,N3308,N3309,N3310,N3311,N3312,N3314,N3315,N3316 
	,N3317,N3318,N3319,N3320,N3321,N3322,N3323,N3324 
	,N3325,N3326,N3327,N3328,N3329,N3330,N3331,N3332 
	,N3333,N3334,N3335,N3336,N3337,N3338,N3339,N3340 
	,N3341,N3342,N3343,N3344,N3345,N3346,N3347,N3349 
	,N3350,N3352,N3353,N3354,N3355,N3356,N3357,N3358 
	,N3359,N3360,N3361,N3362,N3363,N3364,N3365,N3366 
	,N3367,N3368,N3369,N3370,N3371,N3372,N3374,N3375 
	,N3376,N3377,N3378,N3379,N3380,N3381,N3382,N3383 
	,N3384,N3385,N3386,N3387,N3389,N3390,N3391,N3392 
	,N3393,N3394,N3395,N3396,N3397,N3398,N3399,N3400 
	,N3401,N3403,N3404,N3405,N3406,N3407,N3408,N3409 
	,N3410,N3411,N3412,N3413,N3414,N3415,N3416,N3417 
	,N3418,N3419,N3420,N3421,N3422,N3423,N3424,N3425 
	,N3426,N3427,N3429,N3430,N3431,N3433,N3434,N3435 
	,N3436,N3437,N3438,N3439,N3440,N3441,N3442,N3443 
	,N3444,N3445,N3446,N3447,N3448,N3450,N3451,N3452 
	,N3453,N3454,N3455,N3456,N3457,N3458,N3459,N3460 
	,N3461,N3462,N3463,N3464,N3465,N3466,N3467,N3468 
	,N3469,N3470,N3471,N3472,N3473,N3474,N3475,N3476 
	,N3477,N3478,N3479,N3480,N3481,N3482,N3483,N3484 
	,N3485,N3486,N3487,N3489,N3490,N3491,N3492,N3493 
	,N3494,N3495,N3496,N3497,N3498,N3499,N3500,N3501 
	,N3502,N3503,N3504,N3506,N3507,N3508,N3509,N3510 
	,N3511,N3513,N3514,N3515,N3516,N3517,N3518,N3519 
	,N3520,N3521,N3522,N3523,N3524,N3525,N3526,N3527 
	,N3528,N3529,N3530,N3531,N3532,N3533,N3534,N3535 
	,N3536,N3537,N3538,N3539,N3540,N3541,N3542,N3543 
	,N3544,N3546,N3547,N3548,N3550,N3551,N3552,N3553 
	,N3554,N3555,N3556,N3557,N3558,N3559,N3560,N3561 
	,N3562,N3563,N3564,N3565,N3566,N3567,N3568,N3569 
	,N3570,N3572,N3573,N3574,N3575,N3576,N3577,N3578 
	,N3579,N3580,N3581,N3582,N3583,N3584,N3585,N3586 
	,N3587,N3589,N3590,N3591,N3592,N3593,N3594,N3595 
	,N3596,N3597,N3598,N3599,N3600,N3601,N3603,N3604 
	,N3605,N3606,N3607,N3608,N3609,N3610,N3611,N3612 
	,N3613,N3614,N3615,N3616,N3617,N3618,N3619,N3621 
	,N3622,N3623,N3624,N3625,N3626,N3628,N3629,N3630 
	,N3631,N3633,N3634,N3635,N3636,N3637,N3638,N3639 
	,N3640,N3641,N3642,N3643,N3644,N3646,N3647,N3648 
	,N3649,N3650,N3652,N3653,N3654,N3656,N3657,N3658 
	,N3659,N3660,N3661,N3662,N3663,N3664,N3665,N3666 
	,N3667,N3668,N3669,N3670,N3671,N3672,N3673,N3674 
	,N3675,N3676,N3677,N3678,N3679,N3680,N3681,N3682 
	,N3683,N3684,N3685,N3686,N3687,N3689,N3690,N3691 
	,N3692,N3693,N3694,N3695,N3696,N3697,N3698,N3699 
	,N3700,N3701,N3702,N3703,N3704,N3705,N3706,N3707 
	,N3708,N3709,N3710,N3711,N3712,N3714,N3715,N3716 
	,N3717,N3719,N3720,N3721,N3722,N3723,N3724,N3725 
	,N3726,N3727,N3728,N3729,N3730,N3731,N3733,N3734 
	,N3735,N3736,N3737,N3738,N3739,N3740,N3741,N3742 
	,N3743,N3744,N3745,N3746,N3747,N3749,N3750,N3751 
	,N3752,N3753,N3754,N3755,N5360,N5469,N5472,N5473 
	,N5474,N5477,N5480,N5482,N5487,N5489,N5495,N5496 
	,N5497,N5499,N5501,N5502,N5505,N5506,N5507,N5509 
	,N5511,N5520,N5521,N5523,N5526,N5528,N5530,N5536 
	,N5539,N5540,N5542,N5544,N5547,N5552,N5554,N5557 
	,N5634,N5662,N5664,N5666,N5672,N5674,N5679,N5688 
	,N5692,N5758,N5761,N5765,N5766,N5771,N5777,N5781 
	,N5786,N5789,N5815,N5816,N5824,N5825,N5831,N5833 
	,N5834,N5835,N5897,N5904,N5906,N5909,N5942,N5946 
	,N5949,N5957,N5964,N5986,N5994,N6004,N6008,N6025 
	,N6044,N6053,N6055,N6060,N6061,N6063,N6064,N6071 
	,N6073,N6078,N6081,N6082,N6083,N6085,N6087,N6089 
	,N6095,N6097,N6100,N6103,N6106,N6107,N6108,N6110 
	,N6112,N6114,N6117,N6120,N6122,N6123,N6126,N6129 
	,N6132,N6134,N6135,N6138,N6144,N6146,N6148,N6150 
	,N6154,N6157,N6158,N6160,N6162,N6168,N6170,N6173 
	,N6177,N6178,N6181,N6183,N6185,N6191,N6192,N6193 
	,N6196,N6199,N6203,N6205,N6207,N6209,N6210,N6214 
	,N6216,N6218,N6221,N6225,N6226,N6228,N6230,N6232 
	,N6234,N6239,N6242,N6244,N6247,N8426,N8434,N8442 
	,N8450,N8456;
NAND2XL inst_cellmath__17_0_I270 (.Y(N1896), .A(b_exp[0]), .B(b_exp[1]));
AND4XL inst_cellmath__17_0_I10369 (.Y(N1898), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3667 (.Y(N8426), .A(b_exp[7]), .B(b_exp[6]), .C(N1898));
NOR2XL hyperpropagate_4_1_A_I3668 (.Y(inst_cellmath__17), .A(N1896), .B(N8426));
NOR2XL inst_cellmath__19__2__I283 (.Y(N1919), .A(b_man[10]), .B(b_man[9]));
NOR2XL inst_cellmath__19__2__I284 (.Y(N1927), .A(b_man[8]), .B(b_man[7]));
NOR2XL inst_cellmath__19__2__I285 (.Y(N1938), .A(b_man[6]), .B(b_man[5]));
NOR2XL inst_cellmath__19__2__I286 (.Y(N1947), .A(b_man[4]), .B(b_man[3]));
OR4X1 inst_cellmath__19__2__I10370 (.Y(N1932), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
OR4X1 inst_cellmath__19__2__I10371 (.Y(N1941), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 inst_cellmath__19__2__I10372 (.Y(N1951), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4X1 inst_cellmath__19__2__I290 (.Y(N1936), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(N1932));
NAND4XL inst_cellmath__19__2__I292 (.Y(N1930), .A(N1919), .B(N1938), .C(N1927), .D(N1947));
NOR4BX1 inst_cellmath__19__2__I10373 (.Y(inst_cellmath__19), .AN(N1936), .B(N1930), .C(N1941), .D(N1951));
NAND2XL cynw_cm_float_mul_ieee_I295 (.Y(inst_cellmath__21), .A(inst_cellmath__17), .B(inst_cellmath__19));
NOR2XL inst_cellmath__13__1__I296 (.Y(N1981), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL inst_cellmath__13__1__I297 (.Y(N1985), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__13__1__I298 (.Y(N1988), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__13__1__I299 (.Y(N1976), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__13__1__I3663 (.Y(inst_cellmath__13), .A(N1981), .B(N1988), .C(N1985), .D(N1976));
NOR2XL cynw_cm_float_mul_ieee_I303 (.Y(N441), .A(inst_cellmath__13), .B(inst_cellmath__21));
NAND2XL inst_cellmath__10_0_I304 (.Y(N2007), .A(a_exp[0]), .B(a_exp[1]));
AND4XL inst_cellmath__10_0_I10374 (.Y(N2009), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL hyperpropagate_4_1_A_I3669 (.Y(N8434), .A(a_exp[7]), .B(a_exp[6]), .C(N2009));
NOR2XL hyperpropagate_4_1_A_I3670 (.Y(inst_cellmath__10), .A(N2007), .B(N8434));
NOR2XL inst_cellmath__12__0__I317 (.Y(N2030), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__12__0__I318 (.Y(N2038), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__12__0__I319 (.Y(N2049), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__12__0__I320 (.Y(N2058), .A(a_man[4]), .B(a_man[3]));
OR4X1 inst_cellmath__12__0__I10375 (.Y(N2043), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
OR4X1 inst_cellmath__12__0__I10376 (.Y(N2052), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__12__0__I10377 (.Y(N2062), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4X1 inst_cellmath__12__0__I324 (.Y(N2047), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(N2043));
NAND4XL inst_cellmath__12__0__I326 (.Y(N2041), .A(N2030), .B(N2049), .C(N2038), .D(N2058));
NOR4BX1 inst_cellmath__12__0__I10378 (.Y(inst_cellmath__12), .AN(N2047), .B(N2041), .C(N2052), .D(N2062));
NAND2XL cynw_cm_float_mul_ieee_I329 (.Y(inst_cellmath__14), .A(inst_cellmath__10), .B(inst_cellmath__12));
NOR2XL inst_cellmath__20__3__I330 (.Y(N2092), .A(b_exp[0]), .B(b_exp[1]));
NOR2XL inst_cellmath__20__3__I331 (.Y(N2096), .A(b_exp[7]), .B(b_exp[6]));
NOR2XL inst_cellmath__20__3__I332 (.Y(N2099), .A(b_exp[5]), .B(b_exp[4]));
NOR2XL inst_cellmath__20__3__I333 (.Y(N2087), .A(b_exp[3]), .B(b_exp[2]));
NAND4XL inst_cellmath__20__3__I3665 (.Y(inst_cellmath__20), .A(N2092), .B(N2099), .C(N2096), .D(N2087));
NOR2XL cynw_cm_float_mul_ieee_I337 (.Y(N440), .A(inst_cellmath__20), .B(inst_cellmath__14));
NOR2BX1 cynw_cm_float_mul_ieee_I338 (.Y(inst_cellmath__15), .AN(inst_cellmath__10), .B(inst_cellmath__12));
NOR2BX1 cynw_cm_float_mul_ieee_I339 (.Y(inst_cellmath__22), .AN(inst_cellmath__17), .B(inst_cellmath__19));
OR4X1 cynw_cm_float_mul_ieee_I340 (.Y(inst_cellmath__26), .A(inst_cellmath__22), .B(inst_cellmath__15), .C(N441), .D(N440));
XOR2XL cynw_cm_float_mul_ieee_I341 (.Y(inst_cellmath__23), .A(a_sign), .B(b_sign));
NAND2BXL inst_cellmath__41_0_I342 (.Y(N2131), .AN(b_sign), .B(inst_cellmath__22));
MX2XL inst_cellmath__41_0_I343 (.Y(N2136), .A(N2131), .B(a_sign), .S0(inst_cellmath__15));
MX2XL inst_cellmath__41_0_I344 (.Y(x[31]), .A(inst_cellmath__23), .B(N2136), .S0(inst_cellmath__26));
INVXL inst_cellmath__24_0_I345 (.Y(N3529), .A(a_man[0]));
INVXL inst_cellmath__24_0_I346 (.Y(N2268), .A(a_man[1]));
INVXL inst_cellmath__24_0_I347 (.Y(N2624), .A(a_man[2]));
INVXL inst_cellmath__24_0_I348 (.Y(N2988), .A(a_man[3]));
INVXL inst_cellmath__24_0_I349 (.Y(N3334), .A(a_man[4]));
INVXL inst_cellmath__24_0_I350 (.Y(N3675), .A(a_man[5]));
INVXL inst_cellmath__24_0_I351 (.Y(N2417), .A(a_man[6]));
INVXL inst_cellmath__24_0_I352 (.Y(N2779), .A(a_man[7]));
INVXL inst_cellmath__24_0_I353 (.Y(N3131), .A(a_man[8]));
INVXL inst_cellmath__24_0_I354 (.Y(N3473), .A(a_man[9]));
INVXL inst_cellmath__24_0_I355 (.Y(N2212), .A(a_man[10]));
INVXL inst_cellmath__24_0_I356 (.Y(N2566), .A(a_man[11]));
INVXL inst_cellmath__24_0_I357 (.Y(N2924), .A(a_man[12]));
INVXL inst_cellmath__24_0_I358 (.Y(N3276), .A(a_man[13]));
INVXL inst_cellmath__24_0_I359 (.Y(N3616), .A(a_man[14]));
INVXL inst_cellmath__24_0_I360 (.Y(N2352), .A(a_man[15]));
INVXL inst_cellmath__24_0_I361 (.Y(N2716), .A(a_man[16]));
INVXL inst_cellmath__24_0_I362 (.Y(N3076), .A(a_man[17]));
INVXL inst_cellmath__24_0_I363 (.Y(N3415), .A(a_man[18]));
INVXL inst_cellmath__24_0_I364 (.Y(N2152), .A(a_man[19]));
INVXL inst_cellmath__24_0_I365 (.Y(N2504), .A(a_man[20]));
INVXL inst_cellmath__24_0_I366 (.Y(N2862), .A(a_man[21]));
INVXL inst_cellmath__24_0_I367 (.Y(N3217), .A(a_man[22]));
INVXL inst_cellmath__24_0_I368 (.Y(N2357), .A(b_man[0]));
NAND2X1 inst_cellmath__24_0_I369 (.Y(N2721), .A(b_man[1]), .B(N2357));
INVXL inst_cellmath__24_0_I370 (.Y(N3361), .A(b_man[1]));
XNOR2X1 inst_cellmath__24_0_I371 (.Y(N2655), .A(N3529), .B(N3361));
OAI22XL inst_cellmath__24_0_I372 (.Y(N2293), .A0(N2655), .A1(N2357), .B0(N3361), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I373 (.Y(N3364), .A(N2268), .B(N3361));
OA22X1 inst_cellmath__24_0_I374 (.Y(N3701), .A0(N3364), .A1(N2357), .B0(N2655), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I375 (.Y(N2448), .A(N2624), .B(N3361));
OAI22XL inst_cellmath__24_0_I376 (.Y(N3705), .A0(N2448), .A1(N2357), .B0(N3364), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I377 (.Y(N3161), .A(N2988), .B(N3361));
OAI22XL inst_cellmath__24_0_I378 (.Y(N2807), .A0(N3161), .A1(N2357), .B0(N2448), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I379 (.Y(N2239), .A(N3334), .B(N3361));
OAI22XL inst_cellmath__24_0_I380 (.Y(N3504), .A0(N2239), .A1(N2357), .B0(N3161), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I381 (.Y(N2956), .A(N3675), .B(N3361));
OAI22XL inst_cellmath__24_0_I382 (.Y(N2593), .A0(N2956), .A1(N2357), .B0(N2239), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I383 (.Y(N3641), .A(N2417), .B(N3361));
OAI22XL inst_cellmath__24_0_I384 (.Y(N3303), .A0(N3641), .A1(N2357), .B0(N2956), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I385 (.Y(N2746), .A(N2779), .B(N3361));
OAI22XL inst_cellmath__24_0_I386 (.Y(N2382), .A0(N2746), .A1(N2357), .B0(N3641), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I387 (.Y(N3445), .A(N3131), .B(N3361));
OAI22XL inst_cellmath__24_0_I388 (.Y(N3102), .A0(N3445), .A1(N2357), .B0(N2746), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I389 (.Y(N2535), .A(N3473), .B(N3361));
OAI22XL inst_cellmath__24_0_I390 (.Y(N2182), .A0(N2535), .A1(N2357), .B0(N3445), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I391 (.Y(N3247), .A(N2212), .B(N3361));
OAI22XL inst_cellmath__24_0_I392 (.Y(N2892), .A0(N3247), .A1(N2357), .B0(N2535), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I393 (.Y(N2319), .A(N2566), .B(N3361));
OAI22XL inst_cellmath__24_0_I394 (.Y(N3586), .A0(N2319), .A1(N2357), .B0(N3247), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I395 (.Y(N3047), .A(N2924), .B(N3361));
OAI22XL inst_cellmath__24_0_I396 (.Y(N2683), .A0(N3047), .A1(N2357), .B0(N2319), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I397 (.Y(N3731), .A(N3276), .B(N3361));
OAI22XL inst_cellmath__24_0_I398 (.Y(N3386), .A0(N3731), .A1(N2357), .B0(N3047), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I399 (.Y(N2832), .A(N3616), .B(N3361));
OAI22XL inst_cellmath__24_0_I400 (.Y(N2472), .A0(N2832), .A1(N2357), .B0(N3731), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I401 (.Y(N3525), .A(N2352), .B(N3361));
OAI22XL inst_cellmath__24_0_I402 (.Y(N3190), .A0(N3525), .A1(N2357), .B0(N2832), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I403 (.Y(N2620), .A(N2716), .B(N3361));
OAI22XL inst_cellmath__24_0_I404 (.Y(N2264), .A0(N2620), .A1(N2357), .B0(N3525), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I405 (.Y(N3330), .A(N3076), .B(N3361));
OAI22XL inst_cellmath__24_0_I406 (.Y(N2984), .A0(N3330), .A1(N2357), .B0(N2620), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I407 (.Y(N2412), .A(N3415), .B(N3361));
OAI22XL inst_cellmath__24_0_I408 (.Y(N3671), .A0(N2412), .A1(N2357), .B0(N3330), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I409 (.Y(N3127), .A(N2152), .B(N3361));
OAI22XL inst_cellmath__24_0_I410 (.Y(N2776), .A0(N3127), .A1(N2357), .B0(N2412), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I411 (.Y(N2207), .A(N2504), .B(N3361));
OAI22XL inst_cellmath__24_0_I412 (.Y(N3468), .A0(N2207), .A1(N2357), .B0(N3127), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I413 (.Y(N2920), .A(N2862), .B(N3361));
OAI22XL inst_cellmath__24_0_I414 (.Y(N2561), .A0(N2920), .A1(N2357), .B0(N2207), .B1(N2721));
XNOR2X1 inst_cellmath__24_0_I415 (.Y(N3610), .A(N3217), .B(N3361));
OAI22XL inst_cellmath__24_0_I416 (.Y(N3272), .A0(N3610), .A1(N2357), .B0(N2920), .B1(N2721));
INVXL inst_cellmath__24_0_I417 (.Y(N2712), .A(N3361));
OAI22XL inst_cellmath__24_0_I418 (.Y(N2348), .A0(N2712), .A1(N2357), .B0(N3610), .B1(N2721));
MXI2XL inst_cellmath__24_0_I419 (.Y(N3070), .A(N2721), .B(N2357), .S0(N2712));
AOI21XL inst_cellmath__24_0_I420 (.Y(N2859), .A0(N2357), .A1(N2721), .B0(N3361));
XNOR2X1 inst_cellmath__24_0_I421 (.Y(N3014), .A(b_man[2]), .B(b_man[1]));
XOR2XL inst_cellmath__24_0_I422 (.Y(N3662), .A(b_man[3]), .B(b_man[1]));
NAND2X1 inst_cellmath__24_0_I423 (.Y(N3357), .A(N3662), .B(N3014));
INVXL inst_cellmath__24_0_I424 (.Y(N2237), .A(b_man[3]));
NAND2XL inst_cellmath__24_0_I425 (.Y(N3154), .A(b_man[1]), .B(b_man[2]));
AND2XL inst_cellmath__24_0_I426 (.Y(N3495), .A(b_man[3]), .B(N3154));
XNOR2X1 inst_cellmath__24_0_I427 (.Y(N2588), .A(N3529), .B(N2237));
OAI22XL inst_cellmath__24_0_I428 (.Y(N2233), .A0(N2588), .A1(N3014), .B0(N2237), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I429 (.Y(N3298), .A(N2268), .B(N2237));
OAI22XL inst_cellmath__24_0_I430 (.Y(N2948), .A0(N3298), .A1(N3014), .B0(N2588), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I431 (.Y(N2373), .A(N2624), .B(N2237));
OAI22XL inst_cellmath__24_0_I432 (.Y(N3635), .A0(N2373), .A1(N3014), .B0(N3298), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I433 (.Y(N3096), .A(N2988), .B(N2237));
OAI22XL inst_cellmath__24_0_I434 (.Y(N2741), .A0(N3096), .A1(N3014), .B0(N2373), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I435 (.Y(N2176), .A(N3334), .B(N2237));
OAI22XL inst_cellmath__24_0_I436 (.Y(N3439), .A0(N2176), .A1(N3014), .B0(N3096), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I437 (.Y(N2885), .A(N3675), .B(N2237));
OAI22XL inst_cellmath__24_0_I438 (.Y(N2527), .A0(N2885), .A1(N3014), .B0(N2176), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I439 (.Y(N3581), .A(N2417), .B(N2237));
OAI22XL inst_cellmath__24_0_I440 (.Y(N3240), .A0(N3581), .A1(N3014), .B0(N2885), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I441 (.Y(N2674), .A(N2779), .B(N2237));
OAI22XL inst_cellmath__24_0_I442 (.Y(N2314), .A0(N2674), .A1(N3014), .B0(N3581), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I443 (.Y(N3381), .A(N3131), .B(N2237));
OAI22XL inst_cellmath__24_0_I444 (.Y(N3040), .A0(N3381), .A1(N3014), .B0(N2674), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I445 (.Y(N2467), .A(N3473), .B(N2237));
OAI22XL inst_cellmath__24_0_I446 (.Y(N3725), .A0(N2467), .A1(N3014), .B0(N3381), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I447 (.Y(N3182), .A(N2212), .B(N2237));
OAI22XL inst_cellmath__24_0_I448 (.Y(N2822), .A0(N3182), .A1(N3014), .B0(N2467), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I449 (.Y(N2259), .A(N2566), .B(N2237));
OAI22XL inst_cellmath__24_0_I450 (.Y(N3519), .A0(N2259), .A1(N3014), .B0(N3182), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I451 (.Y(N2978), .A(N2924), .B(N2237));
OAI22XL inst_cellmath__24_0_I452 (.Y(N2615), .A0(N2978), .A1(N3014), .B0(N2259), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I453 (.Y(N3665), .A(N3276), .B(N2237));
OAI22XL inst_cellmath__24_0_I454 (.Y(N3324), .A0(N3665), .A1(N3014), .B0(N2978), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I455 (.Y(N2768), .A(N3616), .B(N2237));
OAI22XL inst_cellmath__24_0_I456 (.Y(N2404), .A0(N2768), .A1(N3014), .B0(N3665), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I457 (.Y(N3462), .A(N2352), .B(N2237));
OAI22XL inst_cellmath__24_0_I458 (.Y(N3120), .A0(N3462), .A1(N3014), .B0(N2768), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I459 (.Y(N2555), .A(N2716), .B(N2237));
OAI22XL inst_cellmath__24_0_I460 (.Y(N2201), .A0(N2555), .A1(N3014), .B0(N3462), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I461 (.Y(N3265), .A(N3076), .B(N2237));
OAI22XL inst_cellmath__24_0_I462 (.Y(N2912), .A0(N3265), .A1(N3014), .B0(N2555), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I463 (.Y(N2340), .A(N3415), .B(N2237));
OAI22XL inst_cellmath__24_0_I464 (.Y(N3605), .A0(N2340), .A1(N3014), .B0(N3265), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I465 (.Y(N3065), .A(N2152), .B(N2237));
OAI22XL inst_cellmath__24_0_I466 (.Y(N2704), .A0(N3065), .A1(N3014), .B0(N2340), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I467 (.Y(N3752), .A(N2504), .B(N2237));
OAI22XL inst_cellmath__24_0_I468 (.Y(N3403), .A0(N3752), .A1(N3014), .B0(N3065), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I469 (.Y(N2852), .A(N2862), .B(N2237));
OAI22XL inst_cellmath__24_0_I470 (.Y(N2493), .A0(N2852), .A1(N3014), .B0(N3752), .B1(N3357));
XNOR2X1 inst_cellmath__24_0_I471 (.Y(N3548), .A(N3217), .B(N2237));
OAI22XL inst_cellmath__24_0_I472 (.Y(N3209), .A0(N3548), .A1(N3014), .B0(N2852), .B1(N3357));
INVXL inst_cellmath__24_0_I473 (.Y(N2640), .A(N2237));
OAI22XL inst_cellmath__24_0_I474 (.Y(N2282), .A0(N2640), .A1(N3014), .B0(N3548), .B1(N3357));
MXI2XL inst_cellmath__24_0_I475 (.Y(N3008), .A(N3357), .B(N3014), .S0(N2640));
AOI21XL inst_cellmath__24_0_I476 (.Y(N2796), .A0(N3014), .A1(N3357), .B0(N2237));
XNOR2X1 inst_cellmath__24_0_I477 (.Y(N2941), .A(b_man[4]), .B(b_man[3]));
XOR2XL inst_cellmath__24_0_I478 (.Y(N2881), .A(b_man[5]), .B(b_man[3]));
NAND2X1 inst_cellmath__24_0_I479 (.Y(N3291), .A(N2881), .B(N2941));
INVXL inst_cellmath__24_0_I480 (.Y(N2377), .A(b_man[5]));
NAND2XL inst_cellmath__24_0_I481 (.Y(N3090), .A(b_man[3]), .B(b_man[4]));
AND2XL inst_cellmath__24_0_I482 (.Y(N3430), .A(b_man[5]), .B(N3090));
XNOR2X1 inst_cellmath__24_0_I483 (.Y(N2520), .A(N3529), .B(N2377));
OAI22XL inst_cellmath__24_0_I484 (.Y(N2168), .A0(N2520), .A1(N2941), .B0(N2377), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I485 (.Y(N3234), .A(N2268), .B(N2377));
OAI22XL inst_cellmath__24_0_I486 (.Y(N2877), .A0(N3234), .A1(N2941), .B0(N2520), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I487 (.Y(N2306), .A(N2624), .B(N2377));
OAI22XL inst_cellmath__24_0_I488 (.Y(N3573), .A0(N2306), .A1(N2941), .B0(N3234), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I489 (.Y(N3034), .A(N2988), .B(N2377));
OAI22XL inst_cellmath__24_0_I490 (.Y(N2668), .A0(N3034), .A1(N2941), .B0(N2306), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I491 (.Y(N3716), .A(N3334), .B(N2377));
OAI22XL inst_cellmath__24_0_I492 (.Y(N3375), .A0(N3716), .A1(N2941), .B0(N3034), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I493 (.Y(N2818), .A(N3675), .B(N2377));
OAI22XL inst_cellmath__24_0_I494 (.Y(N2461), .A0(N2818), .A1(N2941), .B0(N3716), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I495 (.Y(N3514), .A(N2417), .B(N2377));
OAI22XL inst_cellmath__24_0_I496 (.Y(N3175), .A0(N3514), .A1(N2941), .B0(N2818), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I497 (.Y(N2608), .A(N2779), .B(N2377));
OAI22XL inst_cellmath__24_0_I498 (.Y(N2255), .A0(N2608), .A1(N2941), .B0(N3514), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I499 (.Y(N3317), .A(N3131), .B(N2377));
OAI22XL inst_cellmath__24_0_I500 (.Y(N2969), .A0(N3317), .A1(N2941), .B0(N2608), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I501 (.Y(N2398), .A(N3473), .B(N2377));
OAI22XL inst_cellmath__24_0_I502 (.Y(N3658), .A0(N2398), .A1(N2941), .B0(N3317), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I503 (.Y(N3114), .A(N2212), .B(N2377));
OAI22XL inst_cellmath__24_0_I504 (.Y(N2760), .A0(N3114), .A1(N2941), .B0(N2398), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I505 (.Y(N2196), .A(N2566), .B(N2377));
OAI22XL inst_cellmath__24_0_I506 (.Y(N3456), .A0(N2196), .A1(N2941), .B0(N3114), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I507 (.Y(N2905), .A(N2924), .B(N2377));
OAI22XL inst_cellmath__24_0_I508 (.Y(N2548), .A0(N2905), .A1(N2941), .B0(N2196), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I509 (.Y(N3598), .A(N3276), .B(N2377));
OAI22XL inst_cellmath__24_0_I510 (.Y(N3259), .A0(N3598), .A1(N2941), .B0(N2905), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I511 (.Y(N2696), .A(N3616), .B(N2377));
OAI22XL inst_cellmath__24_0_I512 (.Y(N2332), .A0(N2696), .A1(N2941), .B0(N3598), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I513 (.Y(N3397), .A(N2352), .B(N2377));
OAI22XL inst_cellmath__24_0_I514 (.Y(N3056), .A0(N3397), .A1(N2941), .B0(N2696), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I515 (.Y(N2485), .A(N2716), .B(N2377));
OAI22XL inst_cellmath__24_0_I516 (.Y(N3745), .A0(N2485), .A1(N2941), .B0(N3397), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I517 (.Y(N3202), .A(N3076), .B(N2377));
OAI22XL inst_cellmath__24_0_I518 (.Y(N2844), .A0(N3202), .A1(N2941), .B0(N2485), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I519 (.Y(N2276), .A(N3415), .B(N2377));
OAI22XL inst_cellmath__24_0_I520 (.Y(N3539), .A0(N2276), .A1(N2941), .B0(N3202), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I521 (.Y(N2997), .A(N2152), .B(N2377));
OAI22XL inst_cellmath__24_0_I522 (.Y(N2633), .A0(N2997), .A1(N2941), .B0(N2276), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I523 (.Y(N3684), .A(N2504), .B(N2377));
OAI22XL inst_cellmath__24_0_I524 (.Y(N3343), .A0(N3684), .A1(N2941), .B0(N2997), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I525 (.Y(N2789), .A(N2862), .B(N2377));
OAI22XL inst_cellmath__24_0_I526 (.Y(N2425), .A0(N2789), .A1(N2941), .B0(N3684), .B1(N3291));
XNOR2X1 inst_cellmath__24_0_I527 (.Y(N3483), .A(N3217), .B(N2377));
OAI22XL inst_cellmath__24_0_I528 (.Y(N3142), .A0(N3483), .A1(N2941), .B0(N2789), .B1(N3291));
INVXL inst_cellmath__24_0_I529 (.Y(N2575), .A(N2377));
OAI22XL inst_cellmath__24_0_I530 (.Y(N2221), .A0(N2575), .A1(N2941), .B0(N3483), .B1(N3291));
MXI2XL inst_cellmath__24_0_I531 (.Y(N2933), .A(N3291), .B(N2941), .S0(N2575));
AOI21XL inst_cellmath__24_0_I532 (.Y(N2726), .A0(N2941), .A1(N3291), .B0(N2377));
XNOR2X1 inst_cellmath__24_0_I533 (.Y(N2871), .A(b_man[6]), .B(b_man[5]));
XOR2XL inst_cellmath__24_0_I534 (.Y(N3691), .A(b_man[7]), .B(b_man[5]));
NAND2X1 inst_cellmath__24_0_I535 (.Y(N3228), .A(N3691), .B(N2871));
INVXL inst_cellmath__24_0_I536 (.Y(N2531), .A(b_man[7]));
NAND2XL inst_cellmath__24_0_I537 (.Y(N3028), .A(b_man[5]), .B(b_man[6]));
AND2XL inst_cellmath__24_0_I538 (.Y(N3369), .A(b_man[7]), .B(N3028));
XNOR2X1 inst_cellmath__24_0_I539 (.Y(N2453), .A(N3529), .B(N2531));
OAI22XL inst_cellmath__24_0_I540 (.Y(N3710), .A0(N2453), .A1(N2871), .B0(N2531), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I541 (.Y(N3168), .A(N2268), .B(N2531));
OAI22XL inst_cellmath__24_0_I542 (.Y(N2813), .A0(N3168), .A1(N2871), .B0(N2453), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I543 (.Y(N2246), .A(N2624), .B(N2531));
OAI22XL inst_cellmath__24_0_I544 (.Y(N3508), .A0(N2246), .A1(N2871), .B0(N3168), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I545 (.Y(N2963), .A(N2988), .B(N2531));
OAI22XL inst_cellmath__24_0_I546 (.Y(N2602), .A0(N2963), .A1(N2871), .B0(N2246), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I547 (.Y(N3648), .A(N3334), .B(N2531));
OAI22XL inst_cellmath__24_0_I548 (.Y(N3310), .A0(N3648), .A1(N2871), .B0(N2963), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I549 (.Y(N2753), .A(N3675), .B(N2531));
OAI22XL inst_cellmath__24_0_I550 (.Y(N2390), .A0(N2753), .A1(N2871), .B0(N3648), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I551 (.Y(N3451), .A(N2417), .B(N2531));
OAI22XL inst_cellmath__24_0_I552 (.Y(N3109), .A0(N3451), .A1(N2871), .B0(N2753), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I553 (.Y(N2542), .A(N2779), .B(N2531));
OAI22XL inst_cellmath__24_0_I554 (.Y(N2188), .A0(N2542), .A1(N2871), .B0(N3451), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I555 (.Y(N3252), .A(N3131), .B(N2531));
OAI22XL inst_cellmath__24_0_I556 (.Y(N2898), .A0(N3252), .A1(N2871), .B0(N2542), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I557 (.Y(N2326), .A(N3473), .B(N2531));
OAI22XL inst_cellmath__24_0_I558 (.Y(N3592), .A0(N2326), .A1(N2871), .B0(N3252), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I559 (.Y(N3052), .A(N2212), .B(N2531));
OAI22XL inst_cellmath__24_0_I560 (.Y(N2689), .A0(N3052), .A1(N2871), .B0(N2326), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I561 (.Y(N3737), .A(N2566), .B(N2531));
OAI22XL inst_cellmath__24_0_I562 (.Y(N3391), .A0(N3737), .A1(N2871), .B0(N3052), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I563 (.Y(N2837), .A(N2924), .B(N2531));
OAI22XL inst_cellmath__24_0_I564 (.Y(N2479), .A0(N2837), .A1(N2871), .B0(N3737), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I565 (.Y(N3531), .A(N3276), .B(N2531));
OAI22XL inst_cellmath__24_0_I566 (.Y(N3194), .A0(N3531), .A1(N2871), .B0(N2837), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I567 (.Y(N2626), .A(N3616), .B(N2531));
OAI22XL inst_cellmath__24_0_I568 (.Y(N2270), .A0(N2626), .A1(N2871), .B0(N3531), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I569 (.Y(N3336), .A(N2352), .B(N2531));
OAI22XL inst_cellmath__24_0_I570 (.Y(N2990), .A0(N3336), .A1(N2871), .B0(N2626), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I571 (.Y(N2419), .A(N2716), .B(N2531));
OAI22XL inst_cellmath__24_0_I572 (.Y(N3677), .A0(N2419), .A1(N2871), .B0(N3336), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I573 (.Y(N3133), .A(N3076), .B(N2531));
OAI22XL inst_cellmath__24_0_I574 (.Y(N2781), .A0(N3133), .A1(N2871), .B0(N2419), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I575 (.Y(N2214), .A(N3415), .B(N2531));
OAI22XL inst_cellmath__24_0_I576 (.Y(N3475), .A0(N2214), .A1(N2871), .B0(N3133), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I577 (.Y(N2925), .A(N2152), .B(N2531));
OAI22XL inst_cellmath__24_0_I578 (.Y(N2568), .A0(N2925), .A1(N2871), .B0(N2214), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I579 (.Y(N3619), .A(N2504), .B(N2531));
OAI22XL inst_cellmath__24_0_I580 (.Y(N3278), .A0(N3619), .A1(N2871), .B0(N2925), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I581 (.Y(N2718), .A(N2862), .B(N2531));
OAI22XL inst_cellmath__24_0_I582 (.Y(N2353), .A0(N2718), .A1(N2871), .B0(N3619), .B1(N3228));
XNOR2X1 inst_cellmath__24_0_I583 (.Y(N3416), .A(N3217), .B(N2531));
OAI22XL inst_cellmath__24_0_I584 (.Y(N3078), .A0(N3416), .A1(N2871), .B0(N2718), .B1(N3228));
INVXL inst_cellmath__24_0_I585 (.Y(N2506), .A(N2531));
OAI22XL inst_cellmath__24_0_I586 (.Y(N2154), .A0(N2506), .A1(N2871), .B0(N3416), .B1(N3228));
MXI2XL inst_cellmath__24_0_I587 (.Y(N2863), .A(N3228), .B(N2871), .S0(N2506));
AOI21XL inst_cellmath__24_0_I588 (.Y(N2653), .A0(N2871), .A1(N3228), .B0(N2531));
XNOR2X1 inst_cellmath__24_0_I589 (.Y(N2805), .A(b_man[8]), .B(b_man[7]));
XOR2XL inst_cellmath__24_0_I590 (.Y(N2911), .A(b_man[9]), .B(b_man[7]));
NAND2X1 inst_cellmath__24_0_I591 (.Y(N3159), .A(N2911), .B(N2805));
INVXL inst_cellmath__24_0_I592 (.Y(N2678), .A(b_man[9]));
NAND2XL inst_cellmath__24_0_I593 (.Y(N2952), .A(b_man[7]), .B(b_man[8]));
AND2XL inst_cellmath__24_0_I594 (.Y(N3301), .A(b_man[9]), .B(N2952));
XNOR2X1 inst_cellmath__24_0_I595 (.Y(N2379), .A(N3529), .B(N2678));
OAI22XL inst_cellmath__24_0_I596 (.Y(N3639), .A0(N2379), .A1(N2805), .B0(N2678), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I597 (.Y(N3101), .A(N2268), .B(N2678));
OAI22XL inst_cellmath__24_0_I598 (.Y(N2744), .A0(N3101), .A1(N2805), .B0(N2379), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I599 (.Y(N2180), .A(N2624), .B(N2678));
OAI22XL inst_cellmath__24_0_I600 (.Y(N3443), .A0(N2180), .A1(N2805), .B0(N3101), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I601 (.Y(N2891), .A(N2988), .B(N2678));
OAI22XL inst_cellmath__24_0_I602 (.Y(N2533), .A0(N2891), .A1(N2805), .B0(N2180), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I603 (.Y(N3585), .A(N3334), .B(N2678));
OAI22XL inst_cellmath__24_0_I604 (.Y(N3245), .A0(N3585), .A1(N2805), .B0(N2891), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I605 (.Y(N2679), .A(N3675), .B(N2678));
OAI22XL inst_cellmath__24_0_I606 (.Y(N2317), .A0(N2679), .A1(N2805), .B0(N3585), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I607 (.Y(N3385), .A(N2417), .B(N2678));
OAI22XL inst_cellmath__24_0_I608 (.Y(N3046), .A0(N3385), .A1(N2805), .B0(N2679), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I609 (.Y(N2471), .A(N2779), .B(N2678));
OAI22XL inst_cellmath__24_0_I610 (.Y(N3729), .A0(N2471), .A1(N2805), .B0(N3385), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I611 (.Y(N3187), .A(N3131), .B(N2678));
OAI22XL inst_cellmath__24_0_I612 (.Y(N2829), .A0(N3187), .A1(N2805), .B0(N2471), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I613 (.Y(N2263), .A(N3473), .B(N2678));
OAI22XL inst_cellmath__24_0_I614 (.Y(N3524), .A0(N2263), .A1(N2805), .B0(N3187), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I615 (.Y(N2983), .A(N2212), .B(N2678));
OAI22XL inst_cellmath__24_0_I616 (.Y(N2618), .A0(N2983), .A1(N2805), .B0(N2263), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I617 (.Y(N3668), .A(N2566), .B(N2678));
OAI22XL inst_cellmath__24_0_I618 (.Y(N3329), .A0(N3668), .A1(N2805), .B0(N2983), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I619 (.Y(N2774), .A(N2924), .B(N2678));
OAI22XL inst_cellmath__24_0_I620 (.Y(N2408), .A0(N2774), .A1(N2805), .B0(N3668), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I621 (.Y(N3466), .A(N3276), .B(N2678));
OAI22XL inst_cellmath__24_0_I622 (.Y(N3125), .A0(N3466), .A1(N2805), .B0(N2774), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I623 (.Y(N2559), .A(N3616), .B(N2678));
OAI22XL inst_cellmath__24_0_I624 (.Y(N2205), .A0(N2559), .A1(N2805), .B0(N3466), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I625 (.Y(N3270), .A(N2352), .B(N2678));
OAI22XL inst_cellmath__24_0_I626 (.Y(N2917), .A0(N3270), .A1(N2805), .B0(N2559), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I627 (.Y(N2346), .A(N2716), .B(N2678));
OAI22XL inst_cellmath__24_0_I628 (.Y(N3608), .A0(N2346), .A1(N2805), .B0(N3270), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I629 (.Y(N3068), .A(N3076), .B(N2678));
OAI22XL inst_cellmath__24_0_I630 (.Y(N2710), .A0(N3068), .A1(N2805), .B0(N2346), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I631 (.Y(N2144), .A(N3415), .B(N2678));
OAI22XL inst_cellmath__24_0_I632 (.Y(N3409), .A0(N2144), .A1(N2805), .B0(N3068), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I633 (.Y(N2857), .A(N2152), .B(N2678));
OAI22XL inst_cellmath__24_0_I634 (.Y(N2498), .A0(N2857), .A1(N2805), .B0(N2144), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I635 (.Y(N3554), .A(N2504), .B(N2678));
OAI22XL inst_cellmath__24_0_I636 (.Y(N3213), .A0(N3554), .A1(N2805), .B0(N2857), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I637 (.Y(N2645), .A(N2862), .B(N2678));
OAI22XL inst_cellmath__24_0_I638 (.Y(N2288), .A0(N2645), .A1(N2805), .B0(N3554), .B1(N3159));
XNOR2X1 inst_cellmath__24_0_I639 (.Y(N3354), .A(N3217), .B(N2678));
OAI22XL inst_cellmath__24_0_I640 (.Y(N3013), .A0(N3354), .A1(N2805), .B0(N2645), .B1(N3159));
INVXL inst_cellmath__24_0_I641 (.Y(N2439), .A(N2678));
OAI22XL inst_cellmath__24_0_I642 (.Y(N3698), .A0(N2439), .A1(N2805), .B0(N3354), .B1(N3159));
MXI2XL inst_cellmath__24_0_I643 (.Y(N2799), .A(N3159), .B(N2805), .S0(N2439));
AOI21XL inst_cellmath__24_0_I644 (.Y(N2586), .A0(N2805), .A1(N3159), .B0(N2678));
XNOR2X1 inst_cellmath__24_0_I645 (.Y(N2737), .A(b_man[10]), .B(b_man[9]));
XOR2XL inst_cellmath__24_0_I646 (.Y(N3720), .A(b_man[11]), .B(b_man[9]));
NAND2X1 inst_cellmath__24_0_I647 (.Y(N3094), .A(N3720), .B(N2737));
INVXL inst_cellmath__24_0_I648 (.Y(N2827), .A(b_man[11]));
NAND2XL inst_cellmath__24_0_I649 (.Y(N2883), .A(b_man[9]), .B(b_man[10]));
AND2XL inst_cellmath__24_0_I650 (.Y(N3236), .A(b_man[11]), .B(N2883));
XNOR2X1 inst_cellmath__24_0_I651 (.Y(N2312), .A(N3529), .B(N2827));
OAI22XL inst_cellmath__24_0_I652 (.Y(N3579), .A0(N2312), .A1(N2737), .B0(N2827), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I653 (.Y(N3038), .A(N2268), .B(N2827));
OAI22XL inst_cellmath__24_0_I654 (.Y(N2671), .A0(N3038), .A1(N2737), .B0(N2312), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I655 (.Y(N3721), .A(N2624), .B(N2827));
OAI22XL inst_cellmath__24_0_I656 (.Y(N3379), .A0(N3721), .A1(N2737), .B0(N3038), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I657 (.Y(N2821), .A(N2988), .B(N2827));
OAI22XL inst_cellmath__24_0_I658 (.Y(N2465), .A0(N2821), .A1(N2737), .B0(N3721), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I659 (.Y(N3518), .A(N3334), .B(N2827));
OAI22XL inst_cellmath__24_0_I660 (.Y(N3178), .A0(N3518), .A1(N2737), .B0(N2821), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I661 (.Y(N2612), .A(N3675), .B(N2827));
OAI22XL inst_cellmath__24_0_I662 (.Y(N2258), .A0(N2612), .A1(N2737), .B0(N3518), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I663 (.Y(N3323), .A(N2417), .B(N2827));
OAI22XL inst_cellmath__24_0_I664 (.Y(N2975), .A0(N3323), .A1(N2737), .B0(N2612), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I665 (.Y(N2403), .A(N2779), .B(N2827));
OAI22XL inst_cellmath__24_0_I666 (.Y(N3661), .A0(N2403), .A1(N2737), .B0(N3323), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I667 (.Y(N3117), .A(N3131), .B(N2827));
OAI22XL inst_cellmath__24_0_I668 (.Y(N2766), .A0(N3117), .A1(N2737), .B0(N2403), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I669 (.Y(N2200), .A(N3473), .B(N2827));
OAI22XL inst_cellmath__24_0_I670 (.Y(N3460), .A0(N2200), .A1(N2737), .B0(N3117), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I671 (.Y(N2910), .A(N2212), .B(N2827));
OAI22XL inst_cellmath__24_0_I672 (.Y(N2552), .A0(N2910), .A1(N2737), .B0(N2200), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I673 (.Y(N3601), .A(N2566), .B(N2827));
OAI22XL inst_cellmath__24_0_I674 (.Y(N3264), .A0(N3601), .A1(N2737), .B0(N2910), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I675 (.Y(N2701), .A(N2924), .B(N2827));
OAI22XL inst_cellmath__24_0_I676 (.Y(N2338), .A0(N2701), .A1(N2737), .B0(N3601), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I677 (.Y(N3401), .A(N3276), .B(N2827));
OAI22XL inst_cellmath__24_0_I678 (.Y(N3061), .A0(N3401), .A1(N2737), .B0(N2701), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I679 (.Y(N2489), .A(N3616), .B(N2827));
OAI22XL inst_cellmath__24_0_I680 (.Y(N3750), .A0(N2489), .A1(N2737), .B0(N3401), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I681 (.Y(N3207), .A(N2352), .B(N2827));
OAI22XL inst_cellmath__24_0_I682 (.Y(N2849), .A0(N3207), .A1(N2737), .B0(N2489), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I683 (.Y(N2280), .A(N2716), .B(N2827));
OAI22XL inst_cellmath__24_0_I684 (.Y(N3544), .A0(N2280), .A1(N2737), .B0(N3207), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I685 (.Y(N3003), .A(N3076), .B(N2827));
OAI22XL inst_cellmath__24_0_I686 (.Y(N2639), .A0(N3003), .A1(N2737), .B0(N2280), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I687 (.Y(N3690), .A(N3415), .B(N2827));
OAI22XL inst_cellmath__24_0_I688 (.Y(N3347), .A0(N3690), .A1(N2737), .B0(N3003), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I689 (.Y(N2794), .A(N2152), .B(N2827));
OAI22XL inst_cellmath__24_0_I690 (.Y(N2429), .A0(N2794), .A1(N2737), .B0(N3690), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I691 (.Y(N3487), .A(N2504), .B(N2827));
OAI22XL inst_cellmath__24_0_I692 (.Y(N3147), .A0(N3487), .A1(N2737), .B0(N2794), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I693 (.Y(N2580), .A(N2862), .B(N2827));
OAI22XL inst_cellmath__24_0_I694 (.Y(N2225), .A0(N2580), .A1(N2737), .B0(N3487), .B1(N3094));
XNOR2X1 inst_cellmath__24_0_I695 (.Y(N3289), .A(N3217), .B(N2827));
OAI22XL inst_cellmath__24_0_I696 (.Y(N2937), .A0(N3289), .A1(N2737), .B0(N2580), .B1(N3094));
INVXL inst_cellmath__24_0_I697 (.Y(N2364), .A(N2827));
OAI22XL inst_cellmath__24_0_I698 (.Y(N3629), .A0(N2364), .A1(N2737), .B0(N3289), .B1(N3094));
MXI2XL inst_cellmath__24_0_I699 (.Y(N2732), .A(N3094), .B(N2737), .S0(N2364));
AOI21XL inst_cellmath__24_0_I700 (.Y(N2518), .A0(N2737), .A1(N3094), .B0(N2827));
XNOR2X1 inst_cellmath__24_0_I701 (.Y(N2664), .A(b_man[12]), .B(b_man[11]));
XOR2XL inst_cellmath__24_0_I702 (.Y(N2942), .A(b_man[13]), .B(b_man[11]));
NAND2X1 inst_cellmath__24_0_I703 (.Y(N3032), .A(N2942), .B(N2664));
INVXL inst_cellmath__24_0_I704 (.Y(N2981), .A(b_man[13]));
NAND2XL inst_cellmath__24_0_I705 (.Y(N2817), .A(b_man[11]), .B(b_man[12]));
AND2XL inst_cellmath__24_0_I706 (.Y(N3172), .A(b_man[13]), .B(N2817));
XNOR2X1 inst_cellmath__24_0_I707 (.Y(N2254), .A(N3529), .B(N2981));
OAI22XL inst_cellmath__24_0_I708 (.Y(N3511), .A0(N2254), .A1(N2664), .B0(N2981), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I709 (.Y(N2966), .A(N2268), .B(N2981));
OAI22XL inst_cellmath__24_0_I710 (.Y(N2604), .A0(N2966), .A1(N2664), .B0(N2254), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I711 (.Y(N3654), .A(N2624), .B(N2981));
OAI22XL inst_cellmath__24_0_I712 (.Y(N3316), .A0(N3654), .A1(N2664), .B0(N2966), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I713 (.Y(N2759), .A(N2988), .B(N2981));
OAI22XL inst_cellmath__24_0_I714 (.Y(N2394), .A0(N2759), .A1(N2664), .B0(N3654), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I715 (.Y(N3453), .A(N3334), .B(N2981));
OAI22XL inst_cellmath__24_0_I716 (.Y(N3111), .A0(N3453), .A1(N2664), .B0(N2759), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I717 (.Y(N2545), .A(N3675), .B(N2981));
OAI22XL inst_cellmath__24_0_I718 (.Y(N2195), .A0(N2545), .A1(N2664), .B0(N3453), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I719 (.Y(N3258), .A(N2417), .B(N2981));
OAI22XL inst_cellmath__24_0_I720 (.Y(N2903), .A0(N3258), .A1(N2664), .B0(N2545), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I721 (.Y(N2330), .A(N2779), .B(N2981));
OAI22XL inst_cellmath__24_0_I722 (.Y(N3595), .A0(N2330), .A1(N2664), .B0(N3258), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I723 (.Y(N3054), .A(N3131), .B(N2981));
OAI22XL inst_cellmath__24_0_I724 (.Y(N2694), .A0(N3054), .A1(N2664), .B0(N2330), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I725 (.Y(N3742), .A(N3473), .B(N2981));
OAI22XL inst_cellmath__24_0_I726 (.Y(N3394), .A0(N3742), .A1(N2664), .B0(N3054), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I727 (.Y(N2841), .A(N2212), .B(N2981));
OAI22XL inst_cellmath__24_0_I728 (.Y(N2482), .A0(N2841), .A1(N2664), .B0(N3742), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I729 (.Y(N3536), .A(N2566), .B(N2981));
OAI22XL inst_cellmath__24_0_I730 (.Y(N3199), .A0(N3536), .A1(N2664), .B0(N2841), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I731 (.Y(N2631), .A(N2924), .B(N2981));
OAI22XL inst_cellmath__24_0_I732 (.Y(N2273), .A0(N2631), .A1(N2664), .B0(N3536), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I733 (.Y(N3340), .A(N3276), .B(N2981));
OAI22XL inst_cellmath__24_0_I734 (.Y(N2994), .A0(N3340), .A1(N2664), .B0(N2631), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I735 (.Y(N2422), .A(N3616), .B(N2981));
OAI22XL inst_cellmath__24_0_I736 (.Y(N3682), .A0(N2422), .A1(N2664), .B0(N3340), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I737 (.Y(N3140), .A(N2352), .B(N2981));
OAI22XL inst_cellmath__24_0_I738 (.Y(N2786), .A0(N3140), .A1(N2664), .B0(N2422), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I739 (.Y(N2218), .A(N2716), .B(N2981));
OAI22XL inst_cellmath__24_0_I740 (.Y(N3479), .A0(N2218), .A1(N2664), .B0(N3140), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I741 (.Y(N2929), .A(N3076), .B(N2981));
OAI22XL inst_cellmath__24_0_I742 (.Y(N2573), .A0(N2929), .A1(N2664), .B0(N2218), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I743 (.Y(N3624), .A(N3415), .B(N2981));
OAI22XL inst_cellmath__24_0_I744 (.Y(N3283), .A0(N3624), .A1(N2664), .B0(N2929), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I745 (.Y(N2723), .A(N2152), .B(N2981));
OAI22XL inst_cellmath__24_0_I746 (.Y(N2359), .A0(N2723), .A1(N2664), .B0(N3624), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I747 (.Y(N3421), .A(N2504), .B(N2981));
OAI22XL inst_cellmath__24_0_I748 (.Y(N3084), .A0(N3421), .A1(N2664), .B0(N2723), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I749 (.Y(N2511), .A(N2862), .B(N2981));
OAI22XL inst_cellmath__24_0_I750 (.Y(N2160), .A0(N2511), .A1(N2664), .B0(N3421), .B1(N3032));
XNOR2X1 inst_cellmath__24_0_I751 (.Y(N3224), .A(N3217), .B(N2981));
OAI22XL inst_cellmath__24_0_I752 (.Y(N2868), .A0(N3224), .A1(N2664), .B0(N2511), .B1(N3032));
INVXL inst_cellmath__24_0_I753 (.Y(N2296), .A(N2981));
OAI22XL inst_cellmath__24_0_I754 (.Y(N3566), .A0(N2296), .A1(N2664), .B0(N3224), .B1(N3032));
MXI2XL inst_cellmath__24_0_I755 (.Y(N2658), .A(N3032), .B(N2664), .S0(N2296));
AOI21XL inst_cellmath__24_0_I756 (.Y(N2451), .A0(N2664), .A1(N3032), .B0(N2981));
XNOR2X1 inst_cellmath__24_0_I757 (.Y(N2598), .A(b_man[14]), .B(b_man[13]));
XOR2XL inst_cellmath__24_0_I758 (.Y(N3751), .A(b_man[15]), .B(b_man[13]));
NAND2X1 inst_cellmath__24_0_I759 (.Y(N2960), .A(N3751), .B(N2598));
INVXL inst_cellmath__24_0_I760 (.Y(N3124), .A(b_man[15]));
NAND2XL inst_cellmath__24_0_I761 (.Y(N2749), .A(b_man[13]), .B(b_man[14]));
AND2XL inst_cellmath__24_0_I762 (.Y(N3105), .A(b_man[15]), .B(N2749));
XNOR2X1 inst_cellmath__24_0_I763 (.Y(N2187), .A(N3529), .B(N3124));
OAI22XL inst_cellmath__24_0_I764 (.Y(N3448), .A0(N2187), .A1(N2598), .B0(N3124), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I765 (.Y(N2895), .A(N2268), .B(N3124));
OAI22XL inst_cellmath__24_0_I766 (.Y(N2537), .A0(N2895), .A1(N2598), .B0(N2187), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I767 (.Y(N3587), .A(N2624), .B(N3124));
OAI22XL inst_cellmath__24_0_I768 (.Y(N3251), .A0(N3587), .A1(N2598), .B0(N2895), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I769 (.Y(N2687), .A(N2988), .B(N3124));
OAI22XL inst_cellmath__24_0_I770 (.Y(N2322), .A0(N2687), .A1(N2598), .B0(N3587), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I771 (.Y(N3387), .A(N3334), .B(N3124));
OAI22XL inst_cellmath__24_0_I772 (.Y(N3048), .A0(N3387), .A1(N2598), .B0(N2687), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I773 (.Y(N2474), .A(N3675), .B(N3124));
OAI22XL inst_cellmath__24_0_I774 (.Y(N3735), .A0(N2474), .A1(N2598), .B0(N3387), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I775 (.Y(N3193), .A(N2417), .B(N3124));
OAI22XL inst_cellmath__24_0_I776 (.Y(N2834), .A0(N3193), .A1(N2598), .B0(N2474), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I777 (.Y(N2266), .A(N2779), .B(N3124));
OAI22XL inst_cellmath__24_0_I778 (.Y(N3526), .A0(N2266), .A1(N2598), .B0(N3193), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I779 (.Y(N2985), .A(N3131), .B(N3124));
OAI22XL inst_cellmath__24_0_I780 (.Y(N2623), .A0(N2985), .A1(N2598), .B0(N2266), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I781 (.Y(N3674), .A(N3473), .B(N3124));
OAI22XL inst_cellmath__24_0_I782 (.Y(N3332), .A0(N3674), .A1(N2598), .B0(N2985), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I783 (.Y(N2778), .A(N2212), .B(N3124));
OAI22XL inst_cellmath__24_0_I784 (.Y(N2414), .A0(N2778), .A1(N2598), .B0(N3674), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I785 (.Y(N3470), .A(N2566), .B(N3124));
OAI22XL inst_cellmath__24_0_I786 (.Y(N3130), .A0(N3470), .A1(N2598), .B0(N2778), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I787 (.Y(N2565), .A(N2924), .B(N3124));
OAI22XL inst_cellmath__24_0_I788 (.Y(N2211), .A0(N2565), .A1(N2598), .B0(N3470), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I789 (.Y(N3274), .A(N3276), .B(N3124));
OAI22XL inst_cellmath__24_0_I790 (.Y(N2921), .A0(N3274), .A1(N2598), .B0(N2565), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I791 (.Y(N2349), .A(N3616), .B(N3124));
OAI22XL inst_cellmath__24_0_I792 (.Y(N3615), .A0(N2349), .A1(N2598), .B0(N3274), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I793 (.Y(N3075), .A(N2352), .B(N3124));
OAI22XL inst_cellmath__24_0_I794 (.Y(N2714), .A0(N3075), .A1(N2598), .B0(N2349), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I795 (.Y(N2149), .A(N2716), .B(N3124));
OAI22XL inst_cellmath__24_0_I796 (.Y(N3412), .A0(N2149), .A1(N2598), .B0(N3075), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I797 (.Y(N2860), .A(N3076), .B(N3124));
OAI22XL inst_cellmath__24_0_I798 (.Y(N2503), .A0(N2860), .A1(N2598), .B0(N2149), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I799 (.Y(N3559), .A(N3415), .B(N3124));
OAI22XL inst_cellmath__24_0_I800 (.Y(N3216), .A0(N3559), .A1(N2598), .B0(N2860), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I801 (.Y(N2650), .A(N2152), .B(N3124));
OAI22XL inst_cellmath__24_0_I802 (.Y(N2290), .A0(N2650), .A1(N2598), .B0(N3559), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I803 (.Y(N3359), .A(N2504), .B(N3124));
OAI22XL inst_cellmath__24_0_I804 (.Y(N3018), .A0(N3359), .A1(N2598), .B0(N2650), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I805 (.Y(N2443), .A(N2862), .B(N3124));
OAI22XL inst_cellmath__24_0_I806 (.Y(N3700), .A0(N2443), .A1(N2598), .B0(N3359), .B1(N2960));
XNOR2X1 inst_cellmath__24_0_I807 (.Y(N3156), .A(N3217), .B(N3124));
OAI22XL inst_cellmath__24_0_I808 (.Y(N2803), .A0(N3156), .A1(N2598), .B0(N2443), .B1(N2960));
INVXL inst_cellmath__24_0_I809 (.Y(N2234), .A(N3124));
OAI22XL inst_cellmath__24_0_I810 (.Y(N3499), .A0(N2234), .A1(N2598), .B0(N3156), .B1(N2960));
MXI2XL inst_cellmath__24_0_I811 (.Y(N2590), .A(N2960), .B(N2598), .S0(N2234));
AOI21XL inst_cellmath__24_0_I812 (.Y(N2376), .A0(N2598), .A1(N2960), .B0(N3124));
XNOR2X1 inst_cellmath__24_0_I813 (.Y(N2529), .A(b_man[16]), .B(b_man[15]));
XOR2XL inst_cellmath__24_0_I814 (.Y(N2973), .A(b_man[17]), .B(b_man[15]));
NAND2X1 inst_cellmath__24_0_I815 (.Y(N2888), .A(N2973), .B(N2529));
INVXL inst_cellmath__24_0_I816 (.Y(N3268), .A(b_man[17]));
NAND2XL inst_cellmath__24_0_I817 (.Y(N2676), .A(b_man[15]), .B(b_man[16]));
AND2XL inst_cellmath__24_0_I818 (.Y(N3043), .A(b_man[17]), .B(N2676));
XNOR2X1 inst_cellmath__24_0_I819 (.Y(N3727), .A(N3529), .B(N3268));
OAI22XL inst_cellmath__24_0_I820 (.Y(N3383), .A0(N3727), .A1(N2529), .B0(N3268), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I821 (.Y(N2826), .A(N2268), .B(N3268));
OAI22XL inst_cellmath__24_0_I822 (.Y(N2469), .A0(N2826), .A1(N2529), .B0(N3727), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I823 (.Y(N3521), .A(N2624), .B(N3268));
OAI22XL inst_cellmath__24_0_I824 (.Y(N3184), .A0(N3521), .A1(N2529), .B0(N2826), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I825 (.Y(N2616), .A(N2988), .B(N3268));
OAI22XL inst_cellmath__24_0_I826 (.Y(N2261), .A0(N2616), .A1(N2529), .B0(N3521), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I827 (.Y(N3327), .A(N3334), .B(N3268));
OAI22XL inst_cellmath__24_0_I828 (.Y(N2979), .A0(N3327), .A1(N2529), .B0(N2616), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I829 (.Y(N2406), .A(N3675), .B(N3268));
OAI22XL inst_cellmath__24_0_I830 (.Y(N3667), .A0(N2406), .A1(N2529), .B0(N3327), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I831 (.Y(N3123), .A(N2417), .B(N3268));
OAI22XL inst_cellmath__24_0_I832 (.Y(N2771), .A0(N3123), .A1(N2529), .B0(N2406), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I833 (.Y(N2203), .A(N2779), .B(N3268));
OAI22XL inst_cellmath__24_0_I834 (.Y(N3463), .A0(N2203), .A1(N2529), .B0(N3123), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I835 (.Y(N2913), .A(N3131), .B(N3268));
OAI22XL inst_cellmath__24_0_I836 (.Y(N2558), .A0(N2913), .A1(N2529), .B0(N2203), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I837 (.Y(N3607), .A(N3473), .B(N3268));
OAI22XL inst_cellmath__24_0_I838 (.Y(N3267), .A0(N3607), .A1(N2529), .B0(N2913), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I839 (.Y(N2706), .A(N2212), .B(N3268));
OAI22XL inst_cellmath__24_0_I840 (.Y(N2341), .A0(N2706), .A1(N2529), .B0(N3607), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I841 (.Y(N3404), .A(N2566), .B(N3268));
OAI22XL inst_cellmath__24_0_I842 (.Y(N3067), .A0(N3404), .A1(N2529), .B0(N2706), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I843 (.Y(N2497), .A(N2924), .B(N3268));
OAI22XL inst_cellmath__24_0_I844 (.Y(N3754), .A0(N2497), .A1(N2529), .B0(N3404), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I845 (.Y(N3211), .A(N3276), .B(N3268));
OAI22XL inst_cellmath__24_0_I846 (.Y(N2853), .A0(N3211), .A1(N2529), .B0(N2497), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I847 (.Y(N2284), .A(N3616), .B(N3268));
OAI22XL inst_cellmath__24_0_I848 (.Y(N3551), .A0(N2284), .A1(N2529), .B0(N3211), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I849 (.Y(N3010), .A(N2352), .B(N3268));
OAI22XL inst_cellmath__24_0_I850 (.Y(N2642), .A0(N3010), .A1(N2529), .B0(N2284), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I851 (.Y(N3693), .A(N2716), .B(N3268));
OAI22XL inst_cellmath__24_0_I852 (.Y(N3350), .A0(N3693), .A1(N2529), .B0(N3010), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I853 (.Y(N2797), .A(N3076), .B(N3268));
OAI22XL inst_cellmath__24_0_I854 (.Y(N2436), .A0(N2797), .A1(N2529), .B0(N3693), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I855 (.Y(N3492), .A(N3415), .B(N3268));
OAI22XL inst_cellmath__24_0_I856 (.Y(N3150), .A0(N3492), .A1(N2529), .B0(N2797), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I857 (.Y(N2583), .A(N2152), .B(N3268));
OAI22XL inst_cellmath__24_0_I858 (.Y(N2228), .A0(N2583), .A1(N2529), .B0(N3492), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I859 (.Y(N3292), .A(N2504), .B(N3268));
OAI22XL inst_cellmath__24_0_I860 (.Y(N2945), .A0(N3292), .A1(N2529), .B0(N2583), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I861 (.Y(N2369), .A(N2862), .B(N3268));
OAI22XL inst_cellmath__24_0_I862 (.Y(N3631), .A0(N2369), .A1(N2529), .B0(N3292), .B1(N2888));
XNOR2X1 inst_cellmath__24_0_I863 (.Y(N3092), .A(N3217), .B(N3268));
OAI22XL inst_cellmath__24_0_I864 (.Y(N2734), .A0(N3092), .A1(N2529), .B0(N2369), .B1(N2888));
INVXL inst_cellmath__24_0_I865 (.Y(N2170), .A(N3268));
OAI22XL inst_cellmath__24_0_I866 (.Y(N3434), .A0(N2170), .A1(N2529), .B0(N3092), .B1(N2888));
MXI2XL inst_cellmath__24_0_I867 (.Y(N2522), .A(N2888), .B(N2529), .S0(N2170));
AOI21XL inst_cellmath__24_0_I868 (.Y(N2309), .A0(N2529), .A1(N2888), .B0(N3268));
XNOR2X1 inst_cellmath__24_0_I869 (.Y(N2463), .A(b_man[18]), .B(b_man[17]));
XOR2XL inst_cellmath__24_0_I870 (.Y(N2169), .A(b_man[19]), .B(b_man[17]));
NAND2X1 inst_cellmath__24_0_I871 (.Y(N2819), .A(N2169), .B(N2463));
INVXL inst_cellmath__24_0_I872 (.Y(N3407), .A(b_man[19]));
NAND2XL inst_cellmath__24_0_I873 (.Y(N2610), .A(b_man[17]), .B(b_man[18]));
AND2XL inst_cellmath__24_0_I874 (.Y(N2971), .A(b_man[19]), .B(N2610));
XNOR2X1 inst_cellmath__24_0_I875 (.Y(N3659), .A(N3529), .B(N3407));
OAI22XL inst_cellmath__24_0_I876 (.Y(N3321), .A0(N3659), .A1(N2463), .B0(N3407), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I877 (.Y(N2763), .A(N2268), .B(N3407));
OAI22XL inst_cellmath__24_0_I878 (.Y(N2400), .A0(N2763), .A1(N2463), .B0(N3659), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I879 (.Y(N3458), .A(N2624), .B(N3407));
OAI22XL inst_cellmath__24_0_I880 (.Y(N3115), .A0(N3458), .A1(N2463), .B0(N2763), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I881 (.Y(N2549), .A(N2988), .B(N3407));
OAI22XL inst_cellmath__24_0_I882 (.Y(N2198), .A0(N2549), .A1(N2463), .B0(N3458), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I883 (.Y(N3261), .A(N3334), .B(N3407));
OAI22XL inst_cellmath__24_0_I884 (.Y(N2907), .A0(N3261), .A1(N2463), .B0(N2549), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I885 (.Y(N2335), .A(N3675), .B(N3407));
OAI22XL inst_cellmath__24_0_I886 (.Y(N3599), .A0(N2335), .A1(N2463), .B0(N3261), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I887 (.Y(N3059), .A(N2417), .B(N3407));
OAI22XL inst_cellmath__24_0_I888 (.Y(N2698), .A0(N3059), .A1(N2463), .B0(N2335), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I889 (.Y(N3747), .A(N2779), .B(N3407));
OAI22XL inst_cellmath__24_0_I890 (.Y(N3399), .A0(N3747), .A1(N2463), .B0(N3059), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I891 (.Y(N2847), .A(N3131), .B(N3407));
OAI22XL inst_cellmath__24_0_I892 (.Y(N2488), .A0(N2847), .A1(N2463), .B0(N3747), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I893 (.Y(N3541), .A(N3473), .B(N3407));
OAI22XL inst_cellmath__24_0_I894 (.Y(N3204), .A0(N3541), .A1(N2463), .B0(N2847), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I895 (.Y(N2635), .A(N2212), .B(N3407));
OAI22XL inst_cellmath__24_0_I896 (.Y(N2278), .A0(N2635), .A1(N2463), .B0(N3541), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I897 (.Y(N3345), .A(N2566), .B(N3407));
OAI22XL inst_cellmath__24_0_I898 (.Y(N3001), .A0(N3345), .A1(N2463), .B0(N2635), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I899 (.Y(N2428), .A(N2924), .B(N3407));
OAI22XL inst_cellmath__24_0_I900 (.Y(N3687), .A0(N2428), .A1(N2463), .B0(N3345), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I901 (.Y(N3144), .A(N3276), .B(N3407));
OAI22XL inst_cellmath__24_0_I902 (.Y(N2791), .A0(N3144), .A1(N2463), .B0(N2428), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I903 (.Y(N2222), .A(N3616), .B(N3407));
OAI22XL inst_cellmath__24_0_I904 (.Y(N3486), .A0(N2222), .A1(N2463), .B0(N3144), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I905 (.Y(N2936), .A(N2352), .B(N3407));
OAI22XL inst_cellmath__24_0_I906 (.Y(N2577), .A0(N2936), .A1(N2463), .B0(N2222), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I907 (.Y(N3626), .A(N2716), .B(N3407));
OAI22XL inst_cellmath__24_0_I908 (.Y(N3286), .A0(N3626), .A1(N2463), .B0(N2936), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I909 (.Y(N2728), .A(N3076), .B(N3407));
OAI22XL inst_cellmath__24_0_I910 (.Y(N2363), .A0(N2728), .A1(N2463), .B0(N3626), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I911 (.Y(N3427), .A(N3415), .B(N3407));
OAI22XL inst_cellmath__24_0_I912 (.Y(N3087), .A0(N3427), .A1(N2463), .B0(N2728), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I913 (.Y(N2516), .A(N2152), .B(N3407));
OAI22XL inst_cellmath__24_0_I914 (.Y(N2163), .A0(N2516), .A1(N2463), .B0(N3427), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I915 (.Y(N3229), .A(N2504), .B(N3407));
OAI22XL inst_cellmath__24_0_I916 (.Y(N2874), .A0(N3229), .A1(N2463), .B0(N2516), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I917 (.Y(N2301), .A(N2862), .B(N3407));
OAI22XL inst_cellmath__24_0_I918 (.Y(N3569), .A0(N2301), .A1(N2463), .B0(N3229), .B1(N2819));
XNOR2X1 inst_cellmath__24_0_I919 (.Y(N3030), .A(N3217), .B(N3407));
OAI22XL inst_cellmath__24_0_I920 (.Y(N2662), .A0(N3030), .A1(N2463), .B0(N2301), .B1(N2819));
INVXL inst_cellmath__24_0_I921 (.Y(N3711), .A(N3407));
OAI22XL inst_cellmath__24_0_I922 (.Y(N3372), .A0(N3711), .A1(N2463), .B0(N3030), .B1(N2819));
MXI2XL inst_cellmath__24_0_I923 (.Y(N2455), .A(N2819), .B(N2463), .S0(N3711));
AOI21XL inst_cellmath__24_0_I924 (.Y(N2250), .A0(N2463), .A1(N2819), .B0(N3407));
XNOR2X1 inst_cellmath__24_0_I925 (.Y(N2392), .A(b_man[20]), .B(b_man[19]));
XOR2XL inst_cellmath__24_0_I926 (.Y(N3007), .A(b_man[21]), .B(b_man[19]));
NAND2X1 inst_cellmath__24_0_I927 (.Y(N2756), .A(N3007), .B(N2392));
INVXL inst_cellmath__24_0_I928 (.Y(N3552), .A(b_man[21]));
NAND2XL inst_cellmath__24_0_I929 (.Y(N2543), .A(b_man[19]), .B(b_man[20]));
AND2XL inst_cellmath__24_0_I930 (.Y(N2901), .A(b_man[21]), .B(N2543));
XNOR2X1 inst_cellmath__24_0_I931 (.Y(N3593), .A(N3529), .B(N3552));
OAI22XL inst_cellmath__24_0_I932 (.Y(N3255), .A0(N3593), .A1(N2392), .B0(N3552), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I933 (.Y(N2691), .A(N2268), .B(N3552));
OAI22XL inst_cellmath__24_0_I934 (.Y(N2328), .A0(N2691), .A1(N2392), .B0(N3593), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I935 (.Y(N3392), .A(N2624), .B(N3552));
OAI22XL inst_cellmath__24_0_I936 (.Y(N3053), .A0(N3392), .A1(N2392), .B0(N2691), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I937 (.Y(N2480), .A(N2988), .B(N3552));
OAI22XL inst_cellmath__24_0_I938 (.Y(N3739), .A0(N2480), .A1(N2392), .B0(N3392), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I939 (.Y(N3196), .A(N3334), .B(N3552));
OAI22XL inst_cellmath__24_0_I940 (.Y(N2839), .A0(N3196), .A1(N2392), .B0(N2480), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I941 (.Y(N2271), .A(N3675), .B(N3552));
OAI22XL inst_cellmath__24_0_I942 (.Y(N3534), .A0(N2271), .A1(N2392), .B0(N3196), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I943 (.Y(N2991), .A(N2417), .B(N3552));
OAI22XL inst_cellmath__24_0_I944 (.Y(N2628), .A0(N2991), .A1(N2392), .B0(N2271), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I945 (.Y(N3679), .A(N2779), .B(N3552));
OAI22XL inst_cellmath__24_0_I946 (.Y(N3337), .A0(N3679), .A1(N2392), .B0(N2991), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I947 (.Y(N2783), .A(N3131), .B(N3552));
OAI22XL inst_cellmath__24_0_I948 (.Y(N2421), .A0(N2783), .A1(N2392), .B0(N3679), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I949 (.Y(N3477), .A(N3473), .B(N3552));
OAI22XL inst_cellmath__24_0_I950 (.Y(N3135), .A0(N3477), .A1(N2392), .B0(N2783), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I951 (.Y(N2570), .A(N2212), .B(N3552));
OAI22XL inst_cellmath__24_0_I952 (.Y(N2216), .A0(N2570), .A1(N2392), .B0(N3477), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I953 (.Y(N3281), .A(N2566), .B(N3552));
OAI22XL inst_cellmath__24_0_I954 (.Y(N2927), .A0(N3281), .A1(N2392), .B0(N2570), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I955 (.Y(N2356), .A(N2924), .B(N3552));
OAI22XL inst_cellmath__24_0_I956 (.Y(N3622), .A0(N2356), .A1(N2392), .B0(N3281), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I957 (.Y(N3081), .A(N3276), .B(N3552));
OAI22XL inst_cellmath__24_0_I958 (.Y(N2720), .A0(N3081), .A1(N2392), .B0(N2356), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I959 (.Y(N2157), .A(N3616), .B(N3552));
OAI22XL inst_cellmath__24_0_I960 (.Y(N3419), .A0(N2157), .A1(N2392), .B0(N3081), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I961 (.Y(N2865), .A(N2352), .B(N3552));
OAI22XL inst_cellmath__24_0_I962 (.Y(N2508), .A0(N2865), .A1(N2392), .B0(N2157), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I963 (.Y(N3562), .A(N2716), .B(N3552));
OAI22XL inst_cellmath__24_0_I964 (.Y(N3222), .A0(N3562), .A1(N2392), .B0(N2865), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I965 (.Y(N2654), .A(N3076), .B(N3552));
OAI22XL inst_cellmath__24_0_I966 (.Y(N2295), .A0(N2654), .A1(N2392), .B0(N3562), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I967 (.Y(N3366), .A(N3415), .B(N3552));
OAI22XL inst_cellmath__24_0_I968 (.Y(N3023), .A0(N3366), .A1(N2392), .B0(N2654), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I969 (.Y(N2447), .A(N2152), .B(N3552));
OAI22XL inst_cellmath__24_0_I970 (.Y(N3704), .A0(N2447), .A1(N2392), .B0(N3366), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I971 (.Y(N3160), .A(N2504), .B(N3552));
OAI22XL inst_cellmath__24_0_I972 (.Y(N2809), .A0(N3160), .A1(N2392), .B0(N2447), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I973 (.Y(N2241), .A(N2862), .B(N3552));
OAI22XL inst_cellmath__24_0_I974 (.Y(N3503), .A0(N2241), .A1(N2392), .B0(N3160), .B1(N2756));
XNOR2X1 inst_cellmath__24_0_I975 (.Y(N2955), .A(N3217), .B(N3552));
OAI22XL inst_cellmath__24_0_I976 (.Y(N2592), .A0(N2955), .A1(N2392), .B0(N2241), .B1(N2756));
INVXL inst_cellmath__24_0_I977 (.Y(N3640), .A(N3552));
OAI22XL inst_cellmath__24_0_I978 (.Y(N3305), .A0(N3640), .A1(N2392), .B0(N2955), .B1(N2756));
MXI2XL inst_cellmath__24_0_I979 (.Y(N2381), .A(N2756), .B(N2392), .S0(N3640));
AOI21XL inst_cellmath__24_0_I980 (.Y(N2183), .A0(N2392), .A1(N2756), .B0(N3552));
XNOR2X1 inst_cellmath__24_0_I981 (.Y(N2318), .A(b_man[22]), .B(b_man[21]));
OR2XL inst_cellmath__24_0_I982 (.Y(N3011), .A(b_man[22]), .B(b_man[21]));
NAND2XL inst_cellmath__24_0_I983 (.Y(N2831), .A(b_man[21]), .B(b_man[22]));
INVXL inst_cellmath__24_0_I984 (.Y(N2775), .A(N3529));
OAI21XL inst_cellmath__24_0_I985 (.Y(N2411), .A0(N2318), .A1(N2775), .B0(N3011));
INVXL inst_cellmath__24_0_I986 (.Y(N3467), .A(N2268));
OAI22XL inst_cellmath__24_0_I987 (.Y(N3128), .A0(N3467), .A1(N2318), .B0(N2775), .B1(N3011));
INVXL inst_cellmath__24_0_I988 (.Y(N2562), .A(N2624));
OAI22XL inst_cellmath__24_0_I989 (.Y(N2206), .A0(N2562), .A1(N2318), .B0(N3467), .B1(N3011));
INVXL inst_cellmath__24_0_I990 (.Y(N3271), .A(N2988));
OAI22XL inst_cellmath__24_0_I991 (.Y(N2919), .A0(N3271), .A1(N2318), .B0(N2562), .B1(N3011));
INVXL inst_cellmath__24_0_I992 (.Y(N2347), .A(N3334));
OAI22XL inst_cellmath__24_0_I993 (.Y(N3611), .A0(N2347), .A1(N2318), .B0(N3271), .B1(N3011));
INVXL inst_cellmath__24_0_I994 (.Y(N3071), .A(N3675));
OAI22XL inst_cellmath__24_0_I995 (.Y(N2711), .A0(N3071), .A1(N2318), .B0(N2347), .B1(N3011));
INVXL inst_cellmath__24_0_I996 (.Y(N2147), .A(N2417));
OAI22XL inst_cellmath__24_0_I997 (.Y(N3410), .A0(N2147), .A1(N2318), .B0(N3071), .B1(N3011));
INVXL inst_cellmath__24_0_I998 (.Y(N2858), .A(N2779));
OAI22XL inst_cellmath__24_0_I999 (.Y(N2500), .A0(N2858), .A1(N2318), .B0(N2147), .B1(N3011));
INVXL inst_cellmath__24_0_I1000 (.Y(N3555), .A(N3131));
OAI22XL inst_cellmath__24_0_I1001 (.Y(N3214), .A0(N3555), .A1(N2318), .B0(N2858), .B1(N3011));
INVXL inst_cellmath__24_0_I1002 (.Y(N2647), .A(N3473));
OAI22XL inst_cellmath__24_0_I1003 (.Y(N2289), .A0(N2647), .A1(N2318), .B0(N3555), .B1(N3011));
INVXL inst_cellmath__24_0_I1004 (.Y(N3356), .A(N2212));
OAI22XL inst_cellmath__24_0_I1005 (.Y(N3015), .A0(N3356), .A1(N2318), .B0(N2647), .B1(N3011));
INVXL inst_cellmath__24_0_I1006 (.Y(N2440), .A(N2566));
OAI22XL inst_cellmath__24_0_I1007 (.Y(N3699), .A0(N2440), .A1(N2318), .B0(N3356), .B1(N3011));
INVXL inst_cellmath__24_0_I1008 (.Y(N3153), .A(N2924));
OAI22XL inst_cellmath__24_0_I1009 (.Y(N2801), .A0(N3153), .A1(N2318), .B0(N2440), .B1(N3011));
INVXL inst_cellmath__24_0_I1010 (.Y(N2232), .A(N3276));
OAI22XL inst_cellmath__24_0_I1011 (.Y(N3496), .A0(N2232), .A1(N2318), .B0(N3153), .B1(N3011));
INVXL inst_cellmath__24_0_I1012 (.Y(N2949), .A(N3616));
OAI22XL inst_cellmath__24_0_I1013 (.Y(N2587), .A0(N2949), .A1(N2318), .B0(N2232), .B1(N3011));
INVXL inst_cellmath__24_0_I1014 (.Y(N3634), .A(N2352));
OAI22XL inst_cellmath__24_0_I1015 (.Y(N3297), .A0(N3634), .A1(N2318), .B0(N2949), .B1(N3011));
INVXL inst_cellmath__24_0_I1016 (.Y(N2740), .A(N2716));
OAI22XL inst_cellmath__24_0_I1017 (.Y(N2374), .A0(N2740), .A1(N2318), .B0(N3634), .B1(N3011));
INVXL inst_cellmath__24_0_I1018 (.Y(N3438), .A(N3076));
OAI22XL inst_cellmath__24_0_I1019 (.Y(N3095), .A0(N3438), .A1(N2318), .B0(N2740), .B1(N3011));
INVXL inst_cellmath__24_0_I1020 (.Y(N2526), .A(N3415));
OAI22XL inst_cellmath__24_0_I1021 (.Y(N2177), .A0(N2526), .A1(N2318), .B0(N3438), .B1(N3011));
INVXL inst_cellmath__24_0_I1022 (.Y(N3241), .A(N2152));
OAI22XL inst_cellmath__24_0_I1023 (.Y(N2884), .A0(N3241), .A1(N2318), .B0(N2526), .B1(N3011));
INVXL inst_cellmath__24_0_I1024 (.Y(N2313), .A(N2504));
OAI22XL inst_cellmath__24_0_I1025 (.Y(N3580), .A0(N2313), .A1(N2318), .B0(N3241), .B1(N3011));
INVXL inst_cellmath__24_0_I1026 (.Y(N3039), .A(N2862));
OAI22XL inst_cellmath__24_0_I1027 (.Y(N2675), .A0(N3039), .A1(N2318), .B0(N2313), .B1(N3011));
INVXL inst_cellmath__24_0_I1028 (.Y(N3726), .A(N3217));
OAI22XL inst_cellmath__24_0_I1029 (.Y(N3380), .A0(N3726), .A1(N2318), .B0(N3039), .B1(N3011));
NOR2XL inst_cellmath__24_0_I1030 (.Y(N2466), .A(N3726), .B(N3011));
INVXL inst_cellmath__24_0_I1031 (.Y(N3183), .A(N2318));
NAND2XL inst_cellmath__24_0_I1032 (.Y(N2977), .A(N2318), .B(N3011));
INVXL inst_cellmath__24_0_I1033 (.Y(N2695), .A(N2859));
INVXL inst_cellmath__24_0_I1034 (.Y(N3057), .A(N2796));
INVXL inst_cellmath__24_0_I1035 (.Y(N3396), .A(N2726));
INVXL inst_cellmath__24_0_I1036 (.Y(N3744), .A(N2653));
INVXL inst_cellmath__24_0_I1037 (.Y(N2487), .A(N2586));
INVXL inst_cellmath__24_0_I1038 (.Y(N2843), .A(N2518));
INVXL inst_cellmath__24_0_I1039 (.Y(N3201), .A(N2451));
INVXL inst_cellmath__24_0_I1040 (.Y(N3540), .A(N2376));
INVXL inst_cellmath__24_0_I1041 (.Y(N2275), .A(N2309));
INVXL inst_cellmath__24_0_I1042 (.Y(N2632), .A(N2250));
INVXL inst_cellmath__24_0_I1043 (.Y(N2998), .A(N2183));
ADDHX1 inst_cellmath__24_0_I1044 (.CO(N3683), .S(N3342), .A(N3495), .B(N3705));
ADDHX1 inst_cellmath__24_0_I1045 (.CO(N2788), .S(N2426), .A(N2807), .B(N2948));
ADDHX1 inst_cellmath__24_0_I1046 (.CO(N3484), .S(N3141), .A(N3430), .B(N3504));
ADDFX1 inst_cellmath__24_0_I1047 (.CO(N2574), .S(N2220), .A(N2168), .B(N3635), .CI(N2788));
ADDHX1 inst_cellmath__24_0_I1048 (.CO(N3285), .S(N2934), .A(N2593), .B(N2741));
ADDFX1 inst_cellmath__24_0_I1049 (.CO(N2362), .S(N3625), .A(N3484), .B(N2877), .CI(N2934));
ADDHX1 inst_cellmath__24_0_I1050 (.CO(N3085), .S(N2725), .A(N3369), .B(N3303));
ADDFX1 inst_cellmath__24_0_I1051 (.CO(N2512), .S(N3148), .A(N3573), .B(N3439), .CI(N3710));
ADDFX1 inst_cellmath__24_0_I1052 (.CO(N2162), .S(N3424), .A(N3285), .B(N2725), .CI(N3148));
ADDHX1 inst_cellmath__24_0_I1053 (.CO(N3227), .S(N2872), .A(N2382), .B(N2527));
ADDFX1 inst_cellmath__24_0_I1054 (.CO(N2661), .S(N2878), .A(N2813), .B(N2668), .CI(N3085));
ADDFX1 inst_cellmath__24_0_I1055 (.CO(N2299), .S(N3567), .A(N2872), .B(N2512), .CI(N2878));
ADDHX1 inst_cellmath__24_0_I1056 (.CO(N3370), .S(N3027), .A(N3301), .B(N3102));
ADDFX1 inst_cellmath__24_0_I1057 (.CO(N2452), .S(N3709), .A(N3375), .B(N3240), .CI(N3508));
ADDFX1 inst_cellmath__24_0_I1058 (.CO(N3507), .S(N2609), .A(N3227), .B(N3639), .CI(N3027));
ADDFX1 inst_cellmath__24_0_I1059 (.CO(N3167), .S(N2814), .A(N2661), .B(N3709), .CI(N2609));
ADDHX1 inst_cellmath__24_0_I1060 (.CO(N2601), .S(N2248), .A(N2182), .B(N2314));
ADDFX1 inst_cellmath__24_0_I1061 (.CO(N3311), .S(N2962), .A(N2602), .B(N2461), .CI(N2744));
ADDFX1 inst_cellmath__24_0_I1062 (.CO(N2754), .S(N2333), .A(N2248), .B(N3370), .CI(N2452));
ADDFX1 inst_cellmath__24_0_I1063 (.CO(N2389), .S(N3647), .A(N3507), .B(N2962), .CI(N2333));
ADDHX1 inst_cellmath__24_0_I1064 (.CO(N3450), .S(N3108), .A(N3236), .B(N2892));
ADDFX1 inst_cellmath__24_0_I1065 (.CO(N2897), .S(N3685), .A(N3175), .B(N3040), .CI(N3310));
ADDFX1 inst_cellmath__24_0_I1066 (.CO(N2541), .S(N2189), .A(N3108), .B(N3311), .CI(N3685));
ADDFX1 inst_cellmath__24_0_I1067 (.CO(N2325), .S(N3425), .A(N3579), .B(N3443), .CI(N2601));
ADDFX1 inst_cellmath__24_0_I1068 (.CO(N3591), .S(N3253), .A(N2189), .B(N2754), .CI(N3425));
ADDHX1 inst_cellmath__24_0_I1069 (.CO(N3051), .S(N2690), .A(N3586), .B(N3725));
ADDFX1 inst_cellmath__24_0_I1070 (.CO(N2478), .S(N3170), .A(N2390), .B(N2255), .CI(N2533));
ADDFX1 inst_cellmath__24_0_I1071 (.CO(N3738), .S(N3390), .A(N2690), .B(N2897), .CI(N3170));
ADDFX1 inst_cellmath__24_0_I1072 (.CO(N3530), .S(N2899), .A(N3450), .B(N2671), .CI(N2325));
ADDFX1 inst_cellmath__24_0_I1073 (.CO(N3195), .S(N2836), .A(N3390), .B(N2541), .CI(N2899));
ADDHX1 inst_cellmath__24_0_I1074 (.CO(N2625), .S(N2269), .A(N3172), .B(N2683));
ADDFX1 inst_cellmath__24_0_I1075 (.CO(N3335), .S(N2989), .A(N2969), .B(N2822), .CI(N3109));
ADDFX1 inst_cellmath__24_0_I1076 (.CO(N2780), .S(N2627), .A(N3379), .B(N3245), .CI(N3511));
ADDFX1 inst_cellmath__24_0_I1077 (.CO(N2420), .S(N3676), .A(N2269), .B(N2478), .CI(N2627));
ADDFX1 inst_cellmath__24_0_I1078 (.CO(N2213), .S(N2355), .A(N2989), .B(N3051), .CI(N3530));
ADDFX1 inst_cellmath__24_0_I1079 (.CO(N3476), .S(N3132), .A(N3738), .B(N3676), .CI(N2355));
ADDHX1 inst_cellmath__24_0_I1080 (.CO(N2926), .S(N2567), .A(N3386), .B(N3519));
ADDFX1 inst_cellmath__24_0_I1081 (.CO(N3618), .S(N3277), .A(N2188), .B(N3658), .CI(N2317));
ADDFX1 inst_cellmath__24_0_I1082 (.CO(N3077), .S(N3703), .A(N2604), .B(N2465), .CI(N2625));
ADDFX1 inst_cellmath__24_0_I1083 (.CO(N2717), .S(N2354), .A(N3335), .B(N3277), .CI(N3703));
ADDFX1 inst_cellmath__24_0_I1084 (.CO(N2505), .S(N3444), .A(N2780), .B(N2567), .CI(N2420));
ADDFX1 inst_cellmath__24_0_I1085 (.CO(N2153), .S(N3418), .A(N2213), .B(N2354), .CI(N3444));
ADDHX1 inst_cellmath__24_0_I1086 (.CO(N3219), .S(N2864), .A(N3105), .B(N2472));
ADDFX1 inst_cellmath__24_0_I1087 (.CO(N2652), .S(N3189), .A(N2760), .B(N2615), .CI(N2898));
ADDFX1 inst_cellmath__24_0_I1088 (.CO(N2292), .S(N3560), .A(N2864), .B(N3618), .CI(N3189));
ADDFX1 inst_cellmath__24_0_I1089 (.CO(N3702), .S(N2918), .A(N3178), .B(N3046), .CI(N3316));
ADDFX1 inst_cellmath__24_0_I1090 (.CO(N3363), .S(N3020), .A(N3448), .B(N2926), .CI(N2918));
ADDFX1 inst_cellmath__24_0_I1091 (.CO(N3158), .S(N2646), .A(N2717), .B(N3077), .CI(N3560));
ADDFX1 inst_cellmath__24_0_I1092 (.CO(N2806), .S(N2444), .A(N3020), .B(N2505), .CI(N2646));
ADDHX1 inst_cellmath__24_0_I1093 (.CO(N2238), .S(N3501), .A(N3190), .B(N3324));
ADDFX1 inst_cellmath__24_0_I1094 (.CO(N3302), .S(N2372), .A(N3592), .B(N3456), .CI(N3729));
ADDFX1 inst_cellmath__24_0_I1095 (.CO(N2951), .S(N2591), .A(N3702), .B(N2652), .CI(N2372));
ADDFX1 inst_cellmath__24_0_I1096 (.CO(N2745), .S(N3724), .A(N2394), .B(N2258), .CI(N2537));
ADDFX1 inst_cellmath__24_0_I1097 (.CO(N2378), .S(N3638), .A(N3219), .B(N3501), .CI(N3724));
ADDFX1 inst_cellmath__24_0_I1098 (.CO(N2181), .S(N3461), .A(N3363), .B(N2292), .CI(N2591));
ADDFX1 inst_cellmath__24_0_I1099 (.CO(N3442), .S(N3100), .A(N3638), .B(N3158), .CI(N3461));
ADDHX1 inst_cellmath__24_0_I1100 (.CO(N2890), .S(N2532), .A(N3043), .B(N2264));
ADDFX1 inst_cellmath__24_0_I1101 (.CO(N3584), .S(N3246), .A(N2548), .B(N2404), .CI(N2689));
ADDFX1 inst_cellmath__24_0_I1102 (.CO(N3045), .S(N3208), .A(N2975), .B(N2829), .CI(N3111));
ADDFX1 inst_cellmath__24_0_I1103 (.CO(N2680), .S(N2316), .A(N2745), .B(N3302), .CI(N3208));
ADDFX1 inst_cellmath__24_0_I1104 (.CO(N2470), .S(N2940), .A(N3383), .B(N3251), .CI(N2238));
ADDFX1 inst_cellmath__24_0_I1105 (.CO(N3730), .S(N3384), .A(N2532), .B(N3246), .CI(N2940));
ADDFX1 inst_cellmath__24_0_I1106 (.CO(N3523), .S(N2667), .A(N2378), .B(N2951), .CI(N2316));
ADDFX1 inst_cellmath__24_0_I1107 (.CO(N3188), .S(N2828), .A(N3384), .B(N2181), .CI(N2667));
ADDHX1 inst_cellmath__24_0_I1108 (.CO(N2619), .S(N2262), .A(N2984), .B(N3120));
ADDFX1 inst_cellmath__24_0_I1109 (.CO(N3328), .S(N2982), .A(N3391), .B(N3259), .CI(N3524));
ADDFX1 inst_cellmath__24_0_I1110 (.CO(N2773), .S(N2397), .A(N2195), .B(N3661), .CI(N2322));
ADDFX1 inst_cellmath__24_0_I1111 (.CO(N2407), .S(N3670), .A(N3045), .B(N3584), .CI(N2397));
ADDFX1 inst_cellmath__24_0_I1112 (.CO(N2204), .S(N3743), .A(N2890), .B(N2469), .CI(N2262));
ADDFX1 inst_cellmath__24_0_I1113 (.CO(N3465), .S(N3126), .A(N2470), .B(N2982), .CI(N3743));
ADDFX1 inst_cellmath__24_0_I1114 (.CO(N3269), .S(N3482), .A(N3730), .B(N2680), .CI(N3670));
ADDFX1 inst_cellmath__24_0_I1115 (.CO(N2916), .S(N2560), .A(N3126), .B(N3523), .CI(N3482));
ADDHX1 inst_cellmath__24_0_I1116 (.CO(N2345), .S(N3609), .A(N2971), .B(N3671));
ADDFX1 inst_cellmath__24_0_I1117 (.CO(N3408), .S(N3226), .A(N2332), .B(N2201), .CI(N2479));
ADDFX1 inst_cellmath__24_0_I1118 (.CO(N3069), .S(N2709), .A(N2773), .B(N3328), .CI(N3226));
ADDFX1 inst_cellmath__24_0_I1119 (.CO(N2856), .S(N2961), .A(N2766), .B(N2618), .CI(N2903));
ADDFX1 inst_cellmath__24_0_I1120 (.CO(N2499), .S(N2143), .A(N2619), .B(N3609), .CI(N2961));
ADDFX1 inst_cellmath__24_0_I1121 (.CO(N2287), .S(N2688), .A(N3184), .B(N3048), .CI(N3321));
ADDFX1 inst_cellmath__24_0_I1122 (.CO(N3553), .S(N3212), .A(N2407), .B(N2204), .CI(N2688));
ADDFX1 inst_cellmath__24_0_I1123 (.CO(N3355), .S(N2418), .A(N3465), .B(N2709), .CI(N2143));
ADDFX1 inst_cellmath__24_0_I1124 (.CO(N3012), .S(N2644), .A(N3269), .B(N3212), .CI(N2418));
ADDHX1 inst_cellmath__24_0_I1125 (.CO(N2438), .S(N3697), .A(N2776), .B(N2912));
ADDFX1 inst_cellmath__24_0_I1126 (.CO(N3493), .S(N2151), .A(N3194), .B(N3056), .CI(N3329));
ADDFX1 inst_cellmath__24_0_I1127 (.CO(N3152), .S(N2800), .A(N2856), .B(N3408), .CI(N2151));
ADDFX1 inst_cellmath__24_0_I1128 (.CO(N2947), .S(N3500), .A(N3595), .B(N3460), .CI(N3735));
ADDFX1 inst_cellmath__24_0_I1129 (.CO(N2585), .S(N2231), .A(N3697), .B(N2287), .CI(N3500));
ADDFX1 inst_cellmath__24_0_I1130 (.CO(N2370), .S(N3244), .A(N2400), .B(N2261), .CI(N2345));
ADDFX1 inst_cellmath__24_0_I1131 (.CO(N3633), .S(N3295), .A(N2499), .B(N3069), .CI(N3244));
ADDFX1 inst_cellmath__24_0_I1132 (.CO(N3436), .S(N2980), .A(N2231), .B(N2800), .CI(N3553));
ADDFX1 inst_cellmath__24_0_I1133 (.CO(N3093), .S(N2739), .A(N3295), .B(N3355), .CI(N2980));
ADDHX1 inst_cellmath__24_0_I1134 (.CO(N2525), .S(N2175), .A(N2901), .B(N3468));
ADDFX1 inst_cellmath__24_0_I1135 (.CO(N3238), .S(N2882), .A(N3745), .B(N3605), .CI(N2270));
ADDFX1 inst_cellmath__24_0_I1136 (.CO(N2673), .S(N2708), .A(N2552), .B(N2408), .CI(N2694));
ADDFX1 inst_cellmath__24_0_I1137 (.CO(N2311), .S(N3578), .A(N2947), .B(N3493), .CI(N2708));
ADDFX1 inst_cellmath__24_0_I1138 (.CO(N3723), .S(N2437), .A(N2979), .B(N2834), .CI(N3115));
ADDFX1 inst_cellmath__24_0_I1139 (.CO(N3378), .S(N3037), .A(N2438), .B(N2175), .CI(N2437));
ADDFX1 inst_cellmath__24_0_I1140 (.CO(N3180), .S(N2173), .A(N2370), .B(N3255), .CI(N2882));
ADDFX1 inst_cellmath__24_0_I1141 (.CO(N2820), .S(N2464), .A(N2585), .B(N3152), .CI(N2173));
ADDFX1 inst_cellmath__24_0_I1142 (.CO(N2614), .S(N3516), .A(N3037), .B(N3578), .CI(N3633));
ADDFX1 inst_cellmath__24_0_I1143 (.CO(N2257), .S(N3517), .A(N3436), .B(N2464), .CI(N3516));
ADDHX1 inst_cellmath__24_0_I1144 (.CO(N3322), .S(N2974), .A(N2561), .B(N2704));
ADDFX1 inst_cellmath__24_0_I1145 (.CO(N2402), .S(N3664), .A(N2990), .B(N2844), .CI(N3125));
ADDFX1 inst_cellmath__24_0_I1146 (.CO(N3459), .S(N3262), .A(N3394), .B(N3264), .CI(N3526));
ADDFX1 inst_cellmath__24_0_I1147 (.CO(N3119), .S(N2765), .A(N2673), .B(N3238), .CI(N3262));
ADDFX1 inst_cellmath__24_0_I1148 (.CO(N2909), .S(N3002), .A(N2198), .B(N3667), .CI(N2328));
ADDFX1 inst_cellmath__24_0_I1149 (.CO(N2554), .S(N2199), .A(N2974), .B(N3723), .CI(N3002));
ADDFX1 inst_cellmath__24_0_I1150 (.CO(N2337), .S(N2730), .A(N3664), .B(N2525), .CI(N2311));
ADDFX1 inst_cellmath__24_0_I1151 (.CO(N3604), .S(N3263), .A(N2199), .B(N2765), .CI(N2730));
ADDFX1 inst_cellmath__24_0_I1152 (.CO(N3400), .S(N2456), .A(N3180), .B(N3378), .CI(N2820));
ADDFX1 inst_cellmath__24_0_I1153 (.CO(N3064), .S(N2700), .A(N2614), .B(N3263), .CI(N2456));
ADDHX1 inst_cellmath__24_0_I1154 (.CO(N2492), .S(N3749), .A(N2831), .B(N2411));
ADDFX1 inst_cellmath__24_0_I1155 (.CO(N3547), .S(N2192), .A(N3272), .B(N3749), .CI(N3403));
ADDFX1 inst_cellmath__24_0_I1156 (.CO(N3206), .S(N2848), .A(N3459), .B(N2402), .CI(N2192));
ADDFX1 inst_cellmath__24_0_I1157 (.CO(N3006), .S(N3535), .A(N3677), .B(N3539), .CI(N2205));
ADDFX1 inst_cellmath__24_0_I1158 (.CO(N2638), .S(N2279), .A(N3322), .B(N2909), .CI(N3535));
ADDFX1 inst_cellmath__24_0_I1159 (.CO(N2432), .S(N3282), .A(N2482), .B(N2338), .CI(N2623));
ADDFX1 inst_cellmath__24_0_I1160 (.CO(N3689), .S(N3346), .A(N2907), .B(N2771), .CI(N3282));
ADDFX1 inst_cellmath__24_0_I1161 (.CO(N3490), .S(N3024), .A(N3119), .B(N3053), .CI(N2554));
ADDFX1 inst_cellmath__24_0_I1162 (.CO(N3146), .S(N2793), .A(N2848), .B(N2337), .CI(N3024));
ADDFX1 inst_cellmath__24_0_I1163 (.CO(N2939), .S(N2748), .A(N3346), .B(N2279), .CI(N3604));
ADDFX1 inst_cellmath__24_0_I1164 (.CO(N2579), .S(N2224), .A(N3400), .B(N2793), .CI(N2748));
ADDHX1 inst_cellmath__24_0_I1165 (.CO(N3628), .S(N3288), .A(N3128), .B(N2492));
ADDFX1 inst_cellmath__24_0_I1166 (.CO(N3088), .S(N2473), .A(N2348), .B(N3288), .CI(N2493));
ADDFX1 inst_cellmath__24_0_I1167 (.CO(N2731), .S(N2366), .A(N3006), .B(N3547), .CI(N2473));
ADDFX1 inst_cellmath__24_0_I1168 (.CO(N2517), .S(N2208), .A(N2781), .B(N2633), .CI(N2917));
ADDFX1 inst_cellmath__24_0_I1169 (.CO(N2166), .S(N3429), .A(N3061), .B(N2432), .CI(N2208));
ADDFX1 inst_cellmath__24_0_I1170 (.CO(N3570), .S(N3556), .A(N3332), .B(N3199), .CI(N3463));
ADDFX1 inst_cellmath__24_0_I1171 (.CO(N3233), .S(N2876), .A(N3739), .B(N3599), .CI(N3556));
ADDFX1 inst_cellmath__24_0_I1172 (.CO(N3031), .S(N3299), .A(N2638), .B(N3206), .CI(N3689));
ADDFX1 inst_cellmath__24_0_I1173 (.CO(N2666), .S(N2304), .A(N2366), .B(N3490), .CI(N3299));
ADDFX1 inst_cellmath__24_0_I1174 (.CO(N2457), .S(N3041), .A(N2876), .B(N3429), .CI(N3146));
ADDFX1 inst_cellmath__24_0_I1175 (.CO(N3714), .S(N3374), .A(N2304), .B(N2939), .CI(N3041));
ADDFX1 inst_cellmath__24_0_I1176 (.CO(N3174), .S(N2816), .A(N2206), .B(N2775), .CI(N3628));
ADDFX1 inst_cellmath__24_0_I1177 (.CO(N2607), .S(N2769), .A(N3070), .B(N3209), .CI(N3343));
ADDFX1 inst_cellmath__24_0_I1178 (.CO(N2253), .S(N3510), .A(N2517), .B(N3088), .CI(N2769));
ADDFX1 inst_cellmath__24_0_I1179 (.CO(N3657), .S(N2494), .A(N3608), .B(N3475), .CI(N3750));
ADDFX1 inst_cellmath__24_0_I1180 (.CO(N3315), .S(N2965), .A(N2816), .B(N3570), .CI(N2494));
ADDFX1 inst_cellmath__24_0_I1181 (.CO(N3113), .S(N2227), .A(N2414), .B(N2273), .CI(N2558));
ADDFX1 inst_cellmath__24_0_I1182 (.CO(N2758), .S(N2393), .A(N2839), .B(N2698), .CI(N2227));
ADDFX1 inst_cellmath__24_0_I1183 (.CO(N2547), .S(N3574), .A(N2166), .B(N2731), .CI(N3233));
ADDFX1 inst_cellmath__24_0_I1184 (.CO(N2194), .S(N3452), .A(N3510), .B(N3031), .CI(N3574));
ADDFX1 inst_cellmath__24_0_I1185 (.CO(N3597), .S(N3319), .A(N2393), .B(N2965), .CI(N2666));
ADDFX1 inst_cellmath__24_0_I1186 (.CO(N3257), .S(N2902), .A(N3452), .B(N2457), .CI(N3319));
INVXL inst_cellmath__24_0_I1187 (.Y(N2845), .A(N3467));
ADDFX1 inst_cellmath__24_0_I1188 (.CO(N2693), .S(N2329), .A(N2282), .B(N2919), .CI(N2845));
ADDFX1 inst_cellmath__24_0_I1189 (.CO(N2840), .S(N2999), .A(N2568), .B(N2425), .CI(N2710));
ADDFX1 inst_cellmath__24_0_I1190 (.CO(N2484), .S(N3741), .A(N3657), .B(N2607), .CI(N2999));
ADDFX1 inst_cellmath__24_0_I1191 (.CO(N2272), .S(N2727), .A(N2994), .B(N2849), .CI(N3130));
ADDFX1 inst_cellmath__24_0_I1192 (.CO(N3538), .S(N3198), .A(N3174), .B(N3113), .CI(N2727));
ADDFX1 inst_cellmath__24_0_I1193 (.CO(N3339), .S(N2454), .A(N3399), .B(N3267), .CI(N3534));
ADDFX1 inst_cellmath__24_0_I1194 (.CO(N2996), .S(N2630), .A(N2329), .B(N2695), .CI(N2454));
ADDFX1 inst_cellmath__24_0_I1195 (.CO(N2785), .S(N2191), .A(N2253), .B(N3315), .CI(N2758));
ADDFX1 inst_cellmath__24_0_I1196 (.CO(N2424), .S(N3681), .A(N2630), .B(N2547), .CI(N2191));
ADDFX1 inst_cellmath__24_0_I1197 (.CO(N2217), .S(N3533), .A(N3198), .B(N3741), .CI(N2194));
ADDFX1 inst_cellmath__24_0_I1198 (.CO(N3481), .S(N3139), .A(N3681), .B(N3597), .CI(N3533));
INVXL inst_cellmath__24_0_I1199 (.Y(N3079), .A(N2562));
ADDFX1 inst_cellmath__24_0_I1200 (.CO(N2931), .S(N2572), .A(N3611), .B(N3467), .CI(N3079));
ADDFX1 inst_cellmath__24_0_I1201 (.CO(N3083), .S(N3220), .A(N3142), .B(N2572), .CI(N3008));
ADDFX1 inst_cellmath__24_0_I1202 (.CO(N2722), .S(N2361), .A(N2840), .B(N2693), .CI(N3220));
ADDFX1 inst_cellmath__24_0_I1203 (.CO(N2510), .S(N2953), .A(N3409), .B(N3278), .CI(N3544));
ADDFX1 inst_cellmath__24_0_I1204 (.CO(N2159), .S(N3423), .A(N3339), .B(N2272), .CI(N2953));
ADDFX1 inst_cellmath__24_0_I1205 (.CO(N3565), .S(N2682), .A(N2211), .B(N3682), .CI(N2341));
ADDFX1 inst_cellmath__24_0_I1206 (.CO(N3223), .S(N2870), .A(N2628), .B(N2488), .CI(N2682));
ADDFX1 inst_cellmath__24_0_I1207 (.CO(N3026), .S(N2410), .A(N2996), .B(N2484), .CI(N3538));
ADDFX1 inst_cellmath__24_0_I1208 (.CO(N2657), .S(N2298), .A(N2361), .B(N2785), .CI(N2410));
ADDFX1 inst_cellmath__24_0_I1209 (.CO(N2450), .S(N2145), .A(N2870), .B(N3423), .CI(N2424));
ADDFX1 inst_cellmath__24_0_I1210 (.CO(N3707), .S(N3368), .A(N2298), .B(N2217), .CI(N2145));
ADDFX1 inst_cellmath__24_0_I1211 (.CO(N3164), .S(N2812), .A(N2562), .B(N3271), .CI(N2711));
ADDFX1 inst_cellmath__24_0_I1212 (.CO(N2597), .S(N3494), .A(N2812), .B(N2931), .CI(N2221));
ADDFX1 inst_cellmath__24_0_I1213 (.CO(N2245), .S(N3506), .A(N2353), .B(N3057), .CI(N3494));
ADDFX1 inst_cellmath__24_0_I1214 (.CO(N3644), .S(N3239), .A(N2639), .B(N2498), .CI(N2786));
ADDFX1 inst_cellmath__24_0_I1215 (.CO(N3309), .S(N2959), .A(N2510), .B(N3083), .CI(N3239));
ADDFX1 inst_cellmath__24_0_I1216 (.CO(N3104), .S(N2976), .A(N3067), .B(N2921), .CI(N3204));
ADDFX1 inst_cellmath__24_0_I1217 (.CO(N2752), .S(N2385), .A(N3337), .B(N3565), .CI(N2976));
ADDFX1 inst_cellmath__24_0_I1218 (.CO(N2540), .S(N2702), .A(N2159), .B(N2722), .CI(N3223));
ADDFX1 inst_cellmath__24_0_I1219 (.CO(N2186), .S(N3447), .A(N2959), .B(N3026), .CI(N2702));
ADDFX1 inst_cellmath__24_0_I1220 (.CO(N3590), .S(N2433), .A(N2385), .B(N3506), .CI(N2657));
ADDFX1 inst_cellmath__24_0_I1221 (.CO(N3250), .S(N2894), .A(N3447), .B(N2450), .CI(N2433));
INVXL inst_cellmath__24_0_I1222 (.Y(N3572), .A(N2347));
ADDFX1 inst_cellmath__24_0_I1223 (.CO(N2686), .S(N2321), .A(N3164), .B(N3410), .CI(N3572));
ADDFX1 inst_cellmath__24_0_I1224 (.CO(N2477), .S(N3734), .A(N3213), .B(N3078), .CI(N2933));
ADDFX1 inst_cellmath__24_0_I1225 (.CO(N3528), .S(N3715), .A(N3479), .B(N3347), .CI(N3615));
ADDFX1 inst_cellmath__24_0_I1226 (.CO(N3192), .S(N2833), .A(N3104), .B(N3644), .CI(N3715));
ADDFX1 inst_cellmath__24_0_I1227 (.CO(N2987), .S(N3455), .A(N2278), .B(N3754), .CI(N2421));
ADDFX1 inst_cellmath__24_0_I1228 (.CO(N2622), .S(N2265), .A(N2321), .B(N2597), .CI(N3455));
ADDFX1 inst_cellmath__24_0_I1229 (.CO(N2416), .S(N3200), .A(N2245), .B(N3734), .CI(N3309));
ADDFX1 inst_cellmath__24_0_I1230 (.CO(N3673), .S(N3331), .A(N2833), .B(N2540), .CI(N3200));
ADDFX1 inst_cellmath__24_0_I1231 (.CO(N3472), .S(N2932), .A(N2265), .B(N2752), .CI(N2186));
ADDFX1 inst_cellmath__24_0_I1232 (.CO(N3129), .S(N2777), .A(N3331), .B(N3590), .CI(N2932));
ADDFX1 inst_cellmath__24_0_I1233 (.CO(N2923), .S(N2660), .A(N2347), .B(N3071), .CI(N2500));
ADDFX1 inst_cellmath__24_0_I1234 (.CO(N2564), .S(N2210), .A(N2288), .B(N2154), .CI(N2660));
ADDFX1 inst_cellmath__24_0_I1235 (.CO(N2351), .S(N2387), .A(N2573), .B(N2429), .CI(N2714));
ADDFX1 inst_cellmath__24_0_I1236 (.CO(N3614), .S(N3273), .A(N3528), .B(N2477), .CI(N2387));
ADDFX1 inst_cellmath__24_0_I1237 (.CO(N3414), .S(N3736), .A(N3001), .B(N2853), .CI(N3135));
ADDFX1 inst_cellmath__24_0_I1238 (.CO(N3074), .S(N2713), .A(N3396), .B(N2987), .CI(N3736));
ADDFX1 inst_cellmath__24_0_I1239 (.CO(N2861), .S(N3474), .A(N2210), .B(N2686), .CI(N3192));
ADDFX1 inst_cellmath__24_0_I1240 (.CO(N2502), .S(N2148), .A(N3273), .B(N2416), .CI(N3474));
ADDFX1 inst_cellmath__24_0_I1241 (.CO(N2291), .S(N3218), .A(N2713), .B(N2622), .CI(N3673));
ADDFX1 inst_cellmath__24_0_I1242 (.CO(N3558), .S(N3215), .A(N2148), .B(N3472), .CI(N3218));
INVXL inst_cellmath__24_0_I1243 (.Y(N2743), .A(N2147));
ADDFX1 inst_cellmath__24_0_I1244 (.CO(N3017), .S(N2649), .A(N2923), .B(N3214), .CI(N2743));
ADDFX1 inst_cellmath__24_0_I1245 (.CO(N3155), .S(N2889), .A(N2863), .B(N3013), .CI(N3147));
ADDFX1 inst_cellmath__24_0_I1246 (.CO(N2804), .S(N2442), .A(N2351), .B(N2564), .CI(N2889));
ADDFX1 inst_cellmath__24_0_I1247 (.CO(N2589), .S(N2617), .A(N3412), .B(N3283), .CI(N3551));
ADDFX1 inst_cellmath__24_0_I1248 (.CO(N2236), .S(N3498), .A(N2649), .B(N3414), .CI(N2617));
ADDFX1 inst_cellmath__24_0_I1249 (.CO(N3636), .S(N2344), .A(N2216), .B(N3687), .CI(N3614));
ADDFX1 inst_cellmath__24_0_I1250 (.CO(N3300), .S(N2950), .A(N2442), .B(N2861), .CI(N2344));
ADDFX1 inst_cellmath__24_0_I1251 (.CO(N3098), .S(N3696), .A(N3498), .B(N3074), .CI(N2502));
ADDFX1 inst_cellmath__24_0_I1252 (.CO(N2742), .S(N2375), .A(N2950), .B(N2291), .CI(N3696));
ADDFX1 inst_cellmath__24_0_I1253 (.CO(N2179), .S(N3441), .A(N2147), .B(N2858), .CI(N2289));
ADDFX1 inst_cellmath__24_0_I1254 (.CO(N3243), .S(N3435), .A(N3698), .B(N3441), .CI(N2225));
ADDFX1 inst_cellmath__24_0_I1255 (.CO(N2887), .S(N2528), .A(N2589), .B(N3155), .CI(N3435));
ADDFX1 inst_cellmath__24_0_I1256 (.CO(N2677), .S(N3177), .A(N2503), .B(N2359), .CI(N2642));
ADDFX1 inst_cellmath__24_0_I1257 (.CO(N2315), .S(N3583), .A(N3017), .B(N3744), .CI(N3177));
ADDFX1 inst_cellmath__24_0_I1258 (.CO(N3728), .S(N2908), .A(N2927), .B(N2791), .CI(N2236));
ADDFX1 inst_cellmath__24_0_I1259 (.CO(N3382), .S(N3042), .A(N2528), .B(N3636), .CI(N2908));
ADDFX1 inst_cellmath__24_0_I1260 (.CO(N3186), .S(N2636), .A(N3583), .B(N2804), .CI(N3300));
ADDFX1 inst_cellmath__24_0_I1261 (.CO(N2825), .S(N2468), .A(N3042), .B(N3098), .CI(N2636));
INVXL inst_cellmath__24_0_I1262 (.Y(N2165), .A(N3555));
ADDFX1 inst_cellmath__24_0_I1263 (.CO(N2260), .S(N3520), .A(N2179), .B(N3015), .CI(N2165));
ADDFX1 inst_cellmath__24_0_I1264 (.CO(N3666), .S(N3326), .A(N3084), .B(N2937), .CI(N2799));
ADDFX1 inst_cellmath__24_0_I1265 (.CO(N3122), .S(N2302), .A(N3350), .B(N3216), .CI(N3486));
ADDFX1 inst_cellmath__24_0_I1266 (.CO(N2770), .S(N2405), .A(N2677), .B(N3243), .CI(N2302));
ADDFX1 inst_cellmath__24_0_I1267 (.CO(N2557), .S(N3653), .A(N3520), .B(N3622), .CI(N3326));
ADDFX1 inst_cellmath__24_0_I1268 (.CO(N2202), .S(N3464), .A(N2315), .B(N2887), .CI(N3653));
ADDFX1 inst_cellmath__24_0_I1269 (.CO(N3606), .S(N3393), .A(N3728), .B(N2405), .CI(N3464));
ADDFX1 inst_cellmath__24_0_I1270 (.CO(N3266), .S(N2915), .A(N3382), .B(N3186), .CI(N3393));
ADDFX1 inst_cellmath__24_0_I1271 (.CO(N3066), .S(N3136), .A(N3555), .B(N2647), .CI(N3699));
ADDFX1 inst_cellmath__24_0_I1272 (.CO(N2705), .S(N2343), .A(N2160), .B(N3629), .CI(N3136));
ADDFX1 inst_cellmath__24_0_I1273 (.CO(N2496), .S(N2867), .A(N2436), .B(N2290), .CI(N2577));
ADDFX1 inst_cellmath__24_0_I1274 (.CO(N3753), .S(N3406), .A(N3122), .B(N3666), .CI(N2867));
ADDFX1 inst_cellmath__24_0_I1275 (.CO(N3550), .S(N2596), .A(N2260), .B(N2720), .CI(N2487));
ADDFX1 inst_cellmath__24_0_I1276 (.CO(N3210), .S(N2855), .A(N2770), .B(N2343), .CI(N2596));
ADDFX1 inst_cellmath__24_0_I1277 (.CO(N3009), .S(N2320), .A(N3406), .B(N2557), .CI(N2202));
ADDFX1 inst_cellmath__24_0_I1278 (.CO(N2641), .S(N2286), .A(N2855), .B(N3606), .CI(N2320));
INVXL inst_cellmath__24_0_I1279 (.Y(N3469), .A(N3356));
ADDFX1 inst_cellmath__24_0_I1280 (.CO(N3692), .S(N3352), .A(N3066), .B(N2801), .CI(N3469));
ADDFX1 inst_cellmath__24_0_I1281 (.CO(N2230), .S(N3612), .A(N2732), .B(N2868), .CI(N3018));
ADDFX1 inst_cellmath__24_0_I1282 (.CO(N3491), .S(N3149), .A(N2496), .B(N2705), .CI(N3612));
ADDFX1 inst_cellmath__24_0_I1283 (.CO(N3293), .S(N3358), .A(N3286), .B(N3150), .CI(N3419));
ADDFX1 inst_cellmath__24_0_I1284 (.CO(N2944), .S(N2582), .A(N3352), .B(N3550), .CI(N3358));
ADDFX1 inst_cellmath__24_0_I1285 (.CO(N2736), .S(N3097), .A(N2582), .B(N3753), .CI(N3149));
ADDFX1 inst_cellmath__24_0_I1286 (.CO(N2368), .S(N3630), .A(N3009), .B(N3210), .CI(N3097));
ADDFX1 inst_cellmath__24_0_I1287 (.CO(N3433), .S(N3091), .A(N3356), .B(N2440), .CI(N3496));
ADDFX1 inst_cellmath__24_0_I1288 (.CO(N2880), .S(N2823), .A(N3566), .B(N3091), .CI(N3700));
ADDFX1 inst_cellmath__24_0_I1289 (.CO(N2521), .S(N2172), .A(N3293), .B(N2230), .CI(N2823));
ADDFX1 inst_cellmath__24_0_I1290 (.CO(N2308), .S(N2556), .A(N2363), .B(N2228), .CI(N2508));
ADDFX1 inst_cellmath__24_0_I1291 (.CO(N3576), .S(N3235), .A(N3692), .B(N2843), .CI(N2556));
ADDFX1 inst_cellmath__24_0_I1292 (.CO(N3377), .S(N2283), .A(N3491), .B(N2944), .CI(N2172));
ADDFX1 inst_cellmath__24_0_I1293 (.CO(N3035), .S(N2670), .A(N3235), .B(N2736), .CI(N2283));
INVXL inst_cellmath__24_0_I1294 (.Y(N3431), .A(N3153));
ADDFX1 inst_cellmath__24_0_I1295 (.CO(N2462), .S(N3719), .A(N3433), .B(N2587), .CI(N3431));
ADDFX1 inst_cellmath__24_0_I1296 (.CO(N2256), .S(N3515), .A(N2945), .B(N2803), .CI(N2658));
ADDFX1 inst_cellmath__24_0_I1297 (.CO(N3320), .S(N3575), .A(N3222), .B(N3087), .CI(N3719));
ADDFX1 inst_cellmath__24_0_I1298 (.CO(N2970), .S(N2611), .A(N2880), .B(N3515), .CI(N3575));
ADDFX1 inst_cellmath__24_0_I1299 (.CO(N2762), .S(N3318), .A(N2521), .B(N2308), .CI(N3576));
ADDFX1 inst_cellmath__24_0_I1300 (.CO(N2399), .S(N3660), .A(N3377), .B(N2611), .CI(N3318));
ADDFX1 inst_cellmath__24_0_I1301 (.CO(N2197), .S(N3058), .A(N3153), .B(N2232), .CI(N3297));
ADDFX1 inst_cellmath__24_0_I1302 (.CO(N3457), .S(N3116), .A(N3631), .B(N3499), .CI(N3058));
ADDFX1 inst_cellmath__24_0_I1303 (.CO(N3260), .S(N2790), .A(N2295), .B(N2163), .CI(N2462));
ADDFX1 inst_cellmath__24_0_I1304 (.CO(N2906), .S(N2551), .A(N3201), .B(N2256), .CI(N2790));
ADDFX1 inst_cellmath__24_0_I1305 (.CO(N2697), .S(N2514), .A(N3116), .B(N3320), .CI(N2970));
ADDFX1 inst_cellmath__24_0_I1306 (.CO(N2334), .S(N3600), .A(N2551), .B(N2762), .CI(N2514));
INVXL inst_cellmath__24_0_I1307 (.Y(N3650), .A(N2949));
ADDFX1 inst_cellmath__24_0_I1308 (.CO(N3398), .S(N3060), .A(N2197), .B(N2374), .CI(N3650));
ADDFX1 inst_cellmath__24_0_I1309 (.CO(N3543), .S(N2190), .A(N2590), .B(N2734), .CI(N2874));
ADDFX1 inst_cellmath__24_0_I1310 (.CO(N3203), .S(N2846), .A(N3260), .B(N3457), .CI(N2190));
ADDFX1 inst_cellmath__24_0_I1311 (.CO(N3000), .S(N3532), .A(N3060), .B(N3023), .CI(N2906));
ADDFX1 inst_cellmath__24_0_I1312 (.CO(N2634), .S(N2277), .A(N2846), .B(N2697), .CI(N3532));
ADDFX1 inst_cellmath__24_0_I1313 (.CO(N3686), .S(N3344), .A(N2949), .B(N3634), .CI(N3095));
ADDFX1 inst_cellmath__24_0_I1314 (.CO(N3143), .S(N3279), .A(N3434), .B(N3344), .CI(N3569));
ADDFX1 inst_cellmath__24_0_I1315 (.CO(N2792), .S(N2427), .A(N3540), .B(N3543), .CI(N3279));
ADDFX1 inst_cellmath__24_0_I1316 (.CO(N2576), .S(N3021), .A(N3398), .B(N3704), .CI(N3203));
ADDFX1 inst_cellmath__24_0_I1317 (.CO(N2223), .S(N3485), .A(N2427), .B(N3000), .CI(N3021));
INVXL inst_cellmath__24_0_I1318 (.Y(N2534), .A(N2740));
ADDFX1 inst_cellmath__24_0_I1319 (.CO(N3287), .S(N2935), .A(N3686), .B(N2177), .CI(N2534));
ADDFX1 inst_cellmath__24_0_I1320 (.CO(N3086), .S(N2729), .A(N2809), .B(N2662), .CI(N2522));
ADDFX1 inst_cellmath__24_0_I1321 (.CO(N2515), .S(N2681), .A(N3143), .B(N2935), .CI(N2729));
ADDFX1 inst_cellmath__24_0_I1322 (.CO(N2164), .S(N3426), .A(N2576), .B(N2792), .CI(N2681));
ADDFX1 inst_cellmath__24_0_I1323 (.CO(N3568), .S(N2409), .A(N2740), .B(N3438), .CI(N2884));
ADDFX1 inst_cellmath__24_0_I1324 (.CO(N3230), .S(N2873), .A(N3503), .B(N3372), .CI(N2409));
ADDFX1 inst_cellmath__24_0_I1325 (.CO(N3029), .S(N2146), .A(N2275), .B(N3287), .CI(N3086));
ADDFX1 inst_cellmath__24_0_I1326 (.CO(N2663), .S(N2300), .A(N2515), .B(N2873), .CI(N2146));
INVXL inst_cellmath__24_0_I1327 (.Y(N3296), .A(N2526));
ADDFX1 inst_cellmath__24_0_I1328 (.CO(N3712), .S(N3371), .A(N3568), .B(N3580), .CI(N3296));
ADDFX1 inst_cellmath__24_0_I1329 (.CO(N2249), .S(N3437), .A(N2455), .B(N2592), .CI(N3371));
ADDFX1 inst_cellmath__24_0_I1330 (.CO(N3509), .S(N3171), .A(N3029), .B(N3230), .CI(N3437));
ADDFX1 inst_cellmath__24_0_I1331 (.CO(N2964), .S(N2603), .A(N2526), .B(N3241), .CI(N2675));
ADDFX1 inst_cellmath__24_0_I1332 (.CO(N2391), .S(N3181), .A(N3305), .B(N2603), .CI(N3712));
ADDFX1 inst_cellmath__24_0_I1333 (.CO(N3652), .S(N3312), .A(N2249), .B(N2632), .CI(N3181));
INVXL inst_cellmath__24_0_I1334 (.Y(N2703), .A(N2313));
ADDFX1 inst_cellmath__24_0_I1335 (.CO(N3110), .S(N2755), .A(N2964), .B(N3380), .CI(N2703));
ADDFX1 inst_cellmath__24_0_I1336 (.CO(N2900), .S(N2544), .A(N2755), .B(N2381), .CI(N2391));
ADDFX1 inst_cellmath__24_0_I1337 (.CO(N2327), .S(N2851), .A(N2313), .B(N3039), .CI(N2466));
ADDFX1 inst_cellmath__24_0_I1338 (.CO(N3594), .S(N3254), .A(N2998), .B(N3110), .CI(N2851));
ADDFX1 inst_cellmath__24_0_I1339 (.CO(N2838), .S(N2481), .A(N3183), .B(N3217), .CI(N2327));
XNOR2X1 inst_cellmath__24_0_I1340 (.Y(N2992), .A(N3217), .B(N2977));
NAND2XL inst_cellmath__24_0_I1341 (.Y(N3678), .A(b_man[1]), .B(N2293));
NOR2XL inst_cellmath__24_0_I1342 (.Y(N2782), .A(N2233), .B(N3342));
NAND2XL inst_cellmath__24_0_I1343 (.Y(N3134), .A(N2233), .B(N3342));
NOR2XL inst_cellmath__24_0_I1344 (.Y(N3478), .A(N3683), .B(N2426));
NAND2XL inst_cellmath__24_0_I1345 (.Y(N2215), .A(N3683), .B(N2426));
NOR2XL inst_cellmath__24_0_I1346 (.Y(N2569), .A(N3141), .B(N2220));
NAND2XL inst_cellmath__24_0_I1347 (.Y(N2928), .A(N3141), .B(N2220));
NOR2XL inst_cellmath__24_0_I1348 (.Y(N3280), .A(N2574), .B(N3625));
NAND2XL inst_cellmath__24_0_I1349 (.Y(N3621), .A(N2574), .B(N3625));
NOR2XL inst_cellmath__24_0_I1350 (.Y(N2358), .A(N2362), .B(N3424));
NAND2XL inst_cellmath__24_0_I1351 (.Y(N2719), .A(N2362), .B(N3424));
NOR2XL inst_cellmath__24_0_I1352 (.Y(N3080), .A(N2162), .B(N3567));
NAND2XL inst_cellmath__24_0_I1353 (.Y(N3420), .A(N2162), .B(N3567));
NOR2XL inst_cellmath__24_0_I1354 (.Y(N2156), .A(N2299), .B(N2814));
NAND2XL inst_cellmath__24_0_I1355 (.Y(N2507), .A(N2299), .B(N2814));
NOR2XL inst_cellmath__24_0_I1356 (.Y(N2866), .A(N3167), .B(N3647));
NAND2XL inst_cellmath__24_0_I1357 (.Y(N3221), .A(N3167), .B(N3647));
NOR2XL inst_cellmath__24_0_I1358 (.Y(N3561), .A(N2389), .B(N3253));
NAND2XL inst_cellmath__24_0_I1359 (.Y(N2294), .A(N2389), .B(N3253));
NOR2XL inst_cellmath__24_0_I1360 (.Y(N2656), .A(N3591), .B(N2836));
NAND2XL inst_cellmath__24_0_I1361 (.Y(N3022), .A(N3591), .B(N2836));
NOR2XL inst_cellmath__24_0_I1362 (.Y(N3365), .A(N3195), .B(N3132));
NAND2XL inst_cellmath__24_0_I1363 (.Y(N3706), .A(N3195), .B(N3132));
NOR2XL inst_cellmath__24_0_I1364 (.Y(N2446), .A(N3476), .B(N3418));
NAND2XL inst_cellmath__24_0_I1365 (.Y(N2808), .A(N3476), .B(N3418));
NOR2XL inst_cellmath__24_0_I1366 (.Y(N3162), .A(N2153), .B(N2444));
NAND2XL inst_cellmath__24_0_I1367 (.Y(N3502), .A(N2153), .B(N2444));
NOR2XL inst_cellmath__24_0_I1368 (.Y(N2240), .A(N2806), .B(N3100));
NAND2XL inst_cellmath__24_0_I1369 (.Y(N2594), .A(N2806), .B(N3100));
NOR2XL inst_cellmath__24_0_I1370 (.Y(N2954), .A(N3442), .B(N2828));
NAND2XL inst_cellmath__24_0_I1371 (.Y(N3304), .A(N3442), .B(N2828));
NOR2XL inst_cellmath__24_0_I1372 (.Y(N3642), .A(N3188), .B(N2560));
NAND2XL inst_cellmath__24_0_I1373 (.Y(N2380), .A(N3188), .B(N2560));
NOR2XL inst_cellmath__24_0_I1374 (.Y(N2747), .A(N2916), .B(N2644));
NAND2XL inst_cellmath__24_0_I1375 (.Y(N3103), .A(N2916), .B(N2644));
NOR2XL inst_cellmath__24_0_I1376 (.Y(N2536), .A(N3701), .B(N3678));
INVXL inst_cellmath__24_0_I1377 (.Y(N3353), .A(N2782));
INVXL inst_cellmath__24_0_I1378 (.Y(N3695), .A(N3134));
OAI21XL inst_cellmath__24_0_I1379 (.Y(N2830), .A0(N3695), .A1(N2536), .B0(N3353));
AOI21XL inst_cellmath__24_0_I1380 (.Y(N2413), .A0(N2215), .A1(N2830), .B0(N3478));
INVXL inst_cellmath__24_0_I1381 (.Y(N2946), .A(N2569));
INVXL inst_cellmath__24_0_I1382 (.Y(N3294), .A(N2928));
OAI21XL inst_cellmath__24_0_I1383 (.Y(N3411), .A0(N3294), .A1(N2413), .B0(N2946));
AOI21XL inst_cellmath__24_0_I1384 (.Y(N2802), .A0(N3621), .A1(N3411), .B0(N3280));
INVXL inst_cellmath__24_0_I1385 (.Y(N3577), .A(N2358));
INVXL inst_cellmath__24_0_I1386 (.Y(N2310), .A(N2719));
OAI21XL inst_cellmath__24_0_I1387 (.Y(N3582), .A0(N2310), .A1(N2802), .B0(N3577));
AOI21XL inst_cellmath__24_0_I1388 (.Y(N2767), .A0(N3420), .A1(N3582), .B0(N3080));
INVXL inst_cellmath__24_0_I1389 (.Y(N2401), .A(N2156));
INVXL inst_cellmath__24_0_I1390 (.Y(N2764), .A(N2507));
OAI21XL inst_cellmath__24_0_I1391 (.Y(N3349), .A0(N2764), .A1(N2767), .B0(N2401));
AOI21XL inst_cellmath__24_0_I1392 (.Y(N2307), .A0(N3221), .A1(N3349), .B0(N2866));
AOI21XL inst_cellmath__24_0_I1393 (.Y(N3717), .A0(N3022), .A1(N3561), .B0(N2656));
NAND2XL inst_cellmath__24_0_I1394 (.Y(N2460), .A(N3022), .B(N2294));
OAI21XL inst_cellmath__24_0_I1395 (.Y(N2486), .A0(N2460), .A1(N2307), .B0(N3717));
AO21XL inst_cellmath__24_0_I1396 (.Y(N3231), .A0(N2808), .A1(N3365), .B0(N2446));
AOI21XL inst_cellmath__24_0_I1397 (.Y(N3169), .A0(N3706), .A1(N2486), .B0(N3365));
AOI31X1 inst_cellmath__24_0_I1398 (.Y(N2247), .A0(N2808), .A1(N3706), .A2(N2486), .B0(N3231));
AOI21XL inst_cellmath__24_0_I1399 (.Y(N3649), .A0(N2594), .A1(N3162), .B0(N2240));
NAND2XL inst_cellmath__24_0_I1400 (.Y(N2388), .A(N2594), .B(N3502));
OAI21XL inst_cellmath__24_0_I1401 (.Y(N3617), .A0(N2388), .A1(N2247), .B0(N3649));
AOI21XL inst_cellmath__24_0_I1402 (.Y(N3417), .A0(N2380), .A1(N2954), .B0(N3642));
NAND2XL inst_cellmath__24_0_I1403 (.Y(N2155), .A(N2380), .B(N3304));
INVXL inst_cellmath__24_0_I1404 (.Y(N2993), .A(N2747));
INVXL inst_cellmath__24_0_I1405 (.Y(N3338), .A(N3103));
INVXL inst_cellmath__24_0_I1406 (.Y(N2784), .A(N3417));
INVXL inst_cellmath__24_0_I1407 (.Y(N3137), .A(N2155));
OAI21XL inst_cellmath__24_0_I1408 (.Y(N3019), .A0(N3338), .A1(N3417), .B0(N2993));
NOR2XL inst_cellmath__24_0_I1409 (.Y(N3362), .A(N3338), .B(N2155));
NOR2BX1 inst_cellmath__24_0_I1410 (.Y(N2209), .AN(N2294), .B(N2307));
NOR2XL inst_cellmath__24_0_I1411 (.Y(N2158), .A(N2209), .B(N3561));
NOR2BX1 inst_cellmath__24_0_I1412 (.Y(N3072), .AN(N3502), .B(N2247));
NOR2XL inst_cellmath__24_0_I1413 (.Y(N3563), .A(N3072), .B(N3162));
AOI21XL inst_cellmath__24_0_I1414 (.Y(N3669), .A0(N3304), .A1(N3617), .B0(N2954));
AOI21XL inst_cellmath__24_0_I1415 (.Y(N2772), .A0(N3137), .A1(N3617), .B0(N2784));
NAND2BXL inst_cellmath__24_0_I1416 (.Y(N2738), .AN(N2782), .B(N3134));
NAND2BXL inst_cellmath__24_0_I1417 (.Y(N2174), .AN(N3478), .B(N2215));
NAND2BXL inst_cellmath__24_0_I1418 (.Y(N3237), .AN(N2569), .B(N2928));
NAND2BXL inst_cellmath__24_0_I1419 (.Y(N2672), .AN(N3280), .B(N3621));
NAND2BXL inst_cellmath__24_0_I1420 (.Y(N3722), .AN(N2358), .B(N2719));
NAND2BXL inst_cellmath__24_0_I1421 (.Y(N3179), .AN(N3080), .B(N3420));
NAND2BXL inst_cellmath__24_0_I1422 (.Y(N2613), .AN(N2156), .B(N2507));
NAND2BXL inst_cellmath__24_0_I1423 (.Y(N3663), .AN(N2866), .B(N3221));
NAND2BXL inst_cellmath__24_0_I1424 (.Y(N3118), .AN(N3561), .B(N2294));
NAND2BXL inst_cellmath__24_0_I1425 (.Y(N2553), .AN(N2656), .B(N3022));
NAND2BXL inst_cellmath__24_0_I1426 (.Y(N3603), .AN(N3365), .B(N3706));
NAND2BXL inst_cellmath__24_0_I1427 (.Y(N3063), .AN(N2446), .B(N2808));
NAND2BXL inst_cellmath__24_0_I1428 (.Y(N2491), .AN(N3162), .B(N3502));
NAND2BXL inst_cellmath__24_0_I1429 (.Y(N3546), .AN(N2240), .B(N2594));
NAND2BXL inst_cellmath__24_0_I1430 (.Y(N3005), .AN(N2954), .B(N3304));
NAND2BXL inst_cellmath__24_0_I1431 (.Y(N2431), .AN(N3642), .B(N2380));
NAND2BXL inst_cellmath__24_0_I1432 (.Y(N3489), .AN(N2747), .B(N3103));
XOR2XL inst_cellmath__24_0_I1433 (.Y(inst_cellmath__24[0]), .A(b_man[1]), .B(N2293));
XOR2XL inst_cellmath__24_0_I1434 (.Y(inst_cellmath__24[1]), .A(N3678), .B(N3701));
XNOR2X1 inst_cellmath__24_0_I1435 (.Y(inst_cellmath__24[2]), .A(N2536), .B(N2738));
XOR2XL inst_cellmath__24_0_I1436 (.Y(inst_cellmath__24[3]), .A(N2830), .B(N2174));
XNOR2X1 inst_cellmath__24_0_I1437 (.Y(inst_cellmath__24[4]), .A(N2413), .B(N3237));
XOR2XL inst_cellmath__24_0_I1438 (.Y(inst_cellmath__24[5]), .A(N3411), .B(N2672));
XNOR2X1 inst_cellmath__24_0_I1439 (.Y(inst_cellmath__24[6]), .A(N2802), .B(N3722));
XOR2XL inst_cellmath__24_0_I1440 (.Y(inst_cellmath__24[7]), .A(N3582), .B(N3179));
XNOR2X1 inst_cellmath__24_0_I1441 (.Y(inst_cellmath__24[8]), .A(N2767), .B(N2613));
XOR2XL inst_cellmath__24_0_I1442 (.Y(inst_cellmath__24[9]), .A(N3349), .B(N3663));
XNOR2X1 inst_cellmath__24_0_I1443 (.Y(inst_cellmath__24[10]), .A(N2307), .B(N3118));
XNOR2X1 inst_cellmath__24_0_I1444 (.Y(inst_cellmath__24[11]), .A(N2158), .B(N2553));
XOR2XL inst_cellmath__24_0_I1445 (.Y(inst_cellmath__24[12]), .A(N2486), .B(N3603));
XNOR2X1 inst_cellmath__24_0_I1446 (.Y(inst_cellmath__24[13]), .A(N3169), .B(N3063));
XNOR2X1 inst_cellmath__24_0_I1447 (.Y(inst_cellmath__24[14]), .A(N2247), .B(N2491));
XNOR2X1 inst_cellmath__24_0_I1448 (.Y(inst_cellmath__24[15]), .A(N3563), .B(N3546));
XOR2XL inst_cellmath__24_0_I1449 (.Y(inst_cellmath__24[16]), .A(N3617), .B(N3005));
XNOR2X1 inst_cellmath__24_0_I1450 (.Y(inst_cellmath__24[17]), .A(N3669), .B(N2431));
XNOR2X1 inst_cellmath__24_0_I1451 (.Y(inst_cellmath__24[18]), .A(N2772), .B(N3489));
AO21XL inst_cellmath__24_0_I1452 (.Y(N2459), .A0(N3362), .A1(N3617), .B0(N3019));
XOR2XL inst_cellmath__24_0_I1453 (.Y(N3513), .A(N3012), .B(N2739));
NOR2XL inst_cellmath__24_0_I1454 (.Y(N2252), .A(N3093), .B(N3517));
XOR2XL inst_cellmath__24_0_I1455 (.Y(N2606), .A(N3093), .B(N3517));
NOR2XL inst_cellmath__24_0_I1456 (.Y(N2968), .A(N2257), .B(N2700));
XOR2XL inst_cellmath__24_0_I1457 (.Y(N3314), .A(N2257), .B(N2700));
NOR2XL inst_cellmath__24_0_I1458 (.Y(N3656), .A(N3064), .B(N2224));
XOR2XL inst_cellmath__24_0_I1459 (.Y(N2396), .A(N3064), .B(N2224));
NOR2XL inst_cellmath__24_0_I1460 (.Y(N2757), .A(N2579), .B(N3374));
XOR2XL inst_cellmath__24_0_I1461 (.Y(N3112), .A(N2579), .B(N3374));
NOR2XL inst_cellmath__24_0_I1462 (.Y(N3454), .A(N3714), .B(N2902));
XOR2XL inst_cellmath__24_0_I1463 (.Y(N2193), .A(N3714), .B(N2902));
NOR2XL inst_cellmath__24_0_I1464 (.Y(N2546), .A(N3257), .B(N3139));
XOR2XL inst_cellmath__24_0_I1465 (.Y(N2904), .A(N3257), .B(N3139));
NOR2XL inst_cellmath__24_0_I1466 (.Y(N3256), .A(N3481), .B(N3368));
XOR2XL inst_cellmath__24_0_I1467 (.Y(N3596), .A(N3481), .B(N3368));
NOR2XL inst_cellmath__24_0_I1468 (.Y(N2331), .A(N3707), .B(N2894));
XOR2XL inst_cellmath__24_0_I1469 (.Y(N2692), .A(N3707), .B(N2894));
NOR2XL inst_cellmath__24_0_I1470 (.Y(N3055), .A(N3250), .B(N2777));
XOR2XL inst_cellmath__24_0_I1471 (.Y(N3395), .A(N3250), .B(N2777));
NOR2XL inst_cellmath__24_0_I1472 (.Y(N3740), .A(N3129), .B(N3215));
XOR2XL inst_cellmath__24_0_I1473 (.Y(N2483), .A(N3129), .B(N3215));
NOR2XL inst_cellmath__24_0_I1474 (.Y(N2842), .A(N3558), .B(N2375));
XOR2XL inst_cellmath__24_0_I1475 (.Y(N3197), .A(N3558), .B(N2375));
NOR2XL inst_cellmath__24_0_I1476 (.Y(N3537), .A(N2742), .B(N2468));
XOR2XL inst_cellmath__24_0_I1477 (.Y(N2274), .A(N2742), .B(N2468));
NOR2XL inst_cellmath__24_0_I1478 (.Y(N2629), .A(N2825), .B(N2915));
XOR2XL inst_cellmath__24_0_I1479 (.Y(N2995), .A(N2825), .B(N2915));
NOR2XL inst_cellmath__24_0_I1480 (.Y(N3341), .A(N3266), .B(N2286));
XOR2XL inst_cellmath__24_0_I1481 (.Y(N3680), .A(N3266), .B(N2286));
NOR2XL inst_cellmath__24_0_I1482 (.Y(N2423), .A(N2641), .B(N3630));
XOR2XL inst_cellmath__24_0_I1483 (.Y(N2787), .A(N2641), .B(N3630));
NOR2XL inst_cellmath__24_0_I1484 (.Y(N3138), .A(N2670), .B(N2368));
XOR2XL inst_cellmath__24_0_I1485 (.Y(N3480), .A(N2670), .B(N2368));
NOR2XL inst_cellmath__24_0_I1486 (.Y(N2219), .A(N3035), .B(N3660));
XOR2XL inst_cellmath__24_0_I1487 (.Y(N2571), .A(N3035), .B(N3660));
NOR2XL inst_cellmath__24_0_I1488 (.Y(N2930), .A(N2399), .B(N3600));
XOR2XL inst_cellmath__24_0_I1489 (.Y(N3284), .A(N2399), .B(N3600));
NOR2XL inst_cellmath__24_0_I1490 (.Y(N3623), .A(N2334), .B(N2277));
XOR2XL inst_cellmath__24_0_I1491 (.Y(N2360), .A(N2334), .B(N2277));
NOR2XL inst_cellmath__24_0_I1492 (.Y(N2724), .A(N2634), .B(N3485));
XOR2XL inst_cellmath__24_0_I1493 (.Y(N3082), .A(N2634), .B(N3485));
NOR2XL inst_cellmath__24_0_I1494 (.Y(N3422), .A(N2223), .B(N3426));
XOR2XL inst_cellmath__24_0_I1495 (.Y(N2161), .A(N2223), .B(N3426));
NOR2XL inst_cellmath__24_0_I1496 (.Y(N2509), .A(N2300), .B(N2164));
XOR2XL inst_cellmath__24_0_I1497 (.Y(N2869), .A(N2300), .B(N2164));
NOR2XL inst_cellmath__24_0_I1498 (.Y(N3225), .A(N2663), .B(N3171));
XOR2XL inst_cellmath__24_0_I1499 (.Y(N3564), .A(N2663), .B(N3171));
NOR2XL inst_cellmath__24_0_I1500 (.Y(N2297), .A(N3509), .B(N3312));
XOR2XL inst_cellmath__24_0_I1501 (.Y(N2659), .A(N3509), .B(N3312));
NOR2XL inst_cellmath__24_0_I1502 (.Y(N3025), .A(N2544), .B(N3652));
XOR2XL inst_cellmath__24_0_I1503 (.Y(N3367), .A(N2544), .B(N3652));
NOR2XL inst_cellmath__24_0_I1504 (.Y(N3708), .A(N3254), .B(N2900));
XOR2XL inst_cellmath__24_0_I1505 (.Y(N2449), .A(N3254), .B(N2900));
NOR2XL inst_cellmath__24_0_I1506 (.Y(N2811), .A(N2481), .B(N3594));
XOR2XL inst_cellmath__24_0_I1507 (.Y(N3166), .A(N2481), .B(N3594));
XNOR2X1 inst_cellmath__24_0_I1508 (.Y(N2244), .A(N2992), .B(N2838));
AOI2BB2X1 inst_cellmath__24_0_I1509 (.Y(N2600), .A0N(N3012), .A1N(N2739), .B0(N2459), .B1(N3513));
AOI21XL inst_cellmath__24_0_I1510 (.Y(N3308), .A0(N3314), .A1(N2252), .B0(N2968));
NAND2XL inst_cellmath__24_0_I1511 (.Y(N3646), .A(N3314), .B(N2606));
AOI21XL inst_cellmath__24_0_I1512 (.Y(N2384), .A0(N3112), .A1(N3656), .B0(N2757));
NAND2XL inst_cellmath__24_0_I1513 (.Y(N2751), .A(N3112), .B(N2396));
AOI21XL inst_cellmath__24_0_I1514 (.Y(N3107), .A0(N2904), .A1(N3454), .B0(N2546));
NAND2XL inst_cellmath__24_0_I1515 (.Y(N3446), .A(N2904), .B(N2193));
AOI21XL inst_cellmath__24_0_I1516 (.Y(N2185), .A0(N2692), .A1(N3256), .B0(N2331));
NAND2XL inst_cellmath__24_0_I1517 (.Y(N2539), .A(N2692), .B(N3596));
AOI21XL inst_cellmath__24_0_I1518 (.Y(N2893), .A0(N2483), .A1(N3055), .B0(N3740));
NAND2XL inst_cellmath__24_0_I1519 (.Y(N3249), .A(N2483), .B(N3395));
AOI21XL inst_cellmath__24_0_I1520 (.Y(N3589), .A0(N2274), .A1(N2842), .B0(N3537));
NAND2XL inst_cellmath__24_0_I1521 (.Y(N2324), .A(N2274), .B(N3197));
AOI21XL inst_cellmath__24_0_I1522 (.Y(N2685), .A0(N3680), .A1(N2629), .B0(N3341));
NAND2XL inst_cellmath__24_0_I1523 (.Y(N3050), .A(N3680), .B(N2995));
AOI21XL inst_cellmath__24_0_I1524 (.Y(N3389), .A0(N3480), .A1(N2423), .B0(N3138));
NAND2XL inst_cellmath__24_0_I1525 (.Y(N3733), .A(N3480), .B(N2787));
AOI21XL inst_cellmath__24_0_I1526 (.Y(N2476), .A0(N3284), .A1(N2219), .B0(N2930));
NAND2XL inst_cellmath__24_0_I1527 (.Y(N2835), .A(N3284), .B(N2571));
AOI21XL inst_cellmath__24_0_I1528 (.Y(N3191), .A0(N3082), .A1(N3623), .B0(N2724));
NAND2XL inst_cellmath__24_0_I1529 (.Y(N3527), .A(N3082), .B(N2360));
AOI21XL inst_cellmath__24_0_I1530 (.Y(N2267), .A0(N2869), .A1(N3422), .B0(N2509));
NAND2XL inst_cellmath__24_0_I1531 (.Y(N2621), .A(N2869), .B(N2161));
AOI21XL inst_cellmath__24_0_I1532 (.Y(N2986), .A0(N2659), .A1(N3225), .B0(N2297));
NAND2XL inst_cellmath__24_0_I1533 (.Y(N3333), .A(N2659), .B(N3564));
AOI21XL inst_cellmath__24_0_I1534 (.Y(N3672), .A0(N2449), .A1(N3025), .B0(N3708));
NAND2XL inst_cellmath__24_0_I1535 (.Y(N2415), .A(N2449), .B(N3367));
OAI21XL inst_cellmath__24_0_I1536 (.Y(N3471), .A0(N3646), .A1(N2600), .B0(N3308));
OAI21XL inst_cellmath__24_0_I1537 (.Y(N2563), .A0(N3446), .A1(N2384), .B0(N3107));
NOR2XL inst_cellmath__24_0_I1538 (.Y(N2922), .A(N3446), .B(N2751));
OAI21XL inst_cellmath__24_0_I1539 (.Y(N3275), .A0(N3249), .A1(N2185), .B0(N2893));
NOR2XL inst_cellmath__24_0_I1540 (.Y(N3613), .A(N3249), .B(N2539));
OAI21XL inst_cellmath__24_0_I1541 (.Y(N2350), .A0(N3050), .A1(N3589), .B0(N2685));
NOR2XL inst_cellmath__24_0_I1542 (.Y(N2715), .A(N3050), .B(N2324));
OAI21XL inst_cellmath__24_0_I1543 (.Y(N3073), .A0(N2835), .A1(N3389), .B0(N2476));
NOR2XL inst_cellmath__24_0_I1544 (.Y(N3413), .A(N2835), .B(N3733));
OAI21XL inst_cellmath__24_0_I1545 (.Y(N2150), .A0(N2621), .A1(N3191), .B0(N2267));
NOR2XL inst_cellmath__24_0_I1546 (.Y(N2501), .A(N2621), .B(N3527));
AOI21XL inst_cellmath__24_0_I1547 (.Y(N3557), .A0(N2922), .A1(N3471), .B0(N2563));
AOI21XL inst_cellmath__24_0_I1548 (.Y(N2651), .A0(N2715), .A1(N3275), .B0(N2350));
NAND2XL inst_cellmath__24_0_I1549 (.Y(N3016), .A(N2715), .B(N3613));
AOI21XL inst_cellmath__24_0_I1550 (.Y(N3360), .A0(N2501), .A1(N3073), .B0(N2150));
OAI21XL inst_cellmath__24_0_I1551 (.Y(N2441), .A0(N3016), .A1(N3557), .B0(N2651));
INVXL inst_cellmath__24_0_I1552 (.Y(N3157), .A(N3613));
INVXL inst_cellmath__24_0_I1553 (.Y(N3497), .A(N3275));
OAI21XL inst_cellmath__24_0_I1554 (.Y(N2235), .A0(N3157), .A1(N3557), .B0(N3497));
INVXL inst_cellmath__24_0_I1555 (.Y(N3163), .A(N2441));
AOI21XL inst_cellmath__24_0_I1556 (.Y(N3637), .A0(N3413), .A1(N2441), .B0(N3073));
INVXL inst_cellmath__24_0_I1557 (.Y(N3099), .A(N3360));
AOI31X1 inst_cellmath__24_0_I1558 (.Y(N3440), .A0(N2501), .A1(N3413), .A2(N2441), .B0(N3099));
INVXL inst_cellmath__24_0_I1559 (.Y(N2530), .A(N2751));
INVXL inst_cellmath__24_0_I1560 (.Y(N2886), .A(N2384));
AOI21XL inst_cellmath__24_0_I1561 (.Y(N3242), .A0(N2530), .A1(N3471), .B0(N2886));
INVXL inst_cellmath__24_0_I1562 (.Y(N2595), .A(N3557));
OAI21XL inst_cellmath__24_0_I1563 (.Y(N3044), .A0(N2539), .A1(N3557), .B0(N2185));
INVXL inst_cellmath__24_0_I1564 (.Y(N2958), .A(N2235));
INVXL inst_cellmath__24_0_I1565 (.Y(N2824), .A(N2324));
INVXL inst_cellmath__24_0_I1566 (.Y(N3185), .A(N3589));
AOI21XL inst_cellmath__24_0_I1567 (.Y(N3522), .A0(N2824), .A1(N2235), .B0(N3185));
INVXL inst_cellmath__24_0_I1568 (.Y(N3306), .A(N3163));
OAI21XL inst_cellmath__24_0_I1569 (.Y(N3325), .A0(N3733), .A1(N3163), .B0(N3389));
INVXL inst_cellmath__24_0_I1570 (.Y(N3643), .A(N3637));
OAI21XL inst_cellmath__24_0_I1571 (.Y(N3121), .A0(N3527), .A1(N3637), .B0(N3191));
INVXL inst_cellmath__24_0_I1572 (.Y(N2383), .A(N3440));
OAI21XL inst_cellmath__24_0_I1573 (.Y(N2914), .A0(N3333), .A1(N3440), .B0(N2986));
OA21X1 inst_cellmath__24_0_I1574 (.Y(N2342), .A0(N2415), .A1(N2986), .B0(N3672));
OAI31X1 inst_cellmath__24_0_I1575 (.Y(N2707), .A0(N2415), .A1(N3333), .A2(N3440), .B0(N2342));
INVXL inst_cellmath__24_0_I1576 (.Y(N3405), .A(N2606));
INVXL inst_cellmath__24_0_I1577 (.Y(N3755), .A(N2252));
OAI21XL inst_cellmath__24_0_I1578 (.Y(N2495), .A0(N3405), .A1(N2600), .B0(N3755));
AOI21XL inst_cellmath__24_0_I1579 (.Y(N2285), .A0(N2396), .A1(N3471), .B0(N3656));
INVXL inst_cellmath__24_0_I1580 (.Y(N3694), .A(N2193));
INVXL inst_cellmath__24_0_I1581 (.Y(N2435), .A(N3454));
OAI21XL inst_cellmath__24_0_I1582 (.Y(N2798), .A0(N3694), .A1(N3242), .B0(N2435));
AOI21XL inst_cellmath__24_0_I1583 (.Y(N2584), .A0(N3596), .A1(N2595), .B0(N3256));
AOI21XL inst_cellmath__24_0_I1584 (.Y(N2367), .A0(N3395), .A1(N3044), .B0(N3055));
INVXL inst_cellmath__24_0_I1585 (.Y(N2171), .A(N3197));
INVXL inst_cellmath__24_0_I1586 (.Y(N2524), .A(N2842));
OAI21XL inst_cellmath__24_0_I1587 (.Y(N2879), .A0(N2171), .A1(N2958), .B0(N2524));
INVXL inst_cellmath__24_0_I1588 (.Y(N2669), .A(N2995));
INVXL inst_cellmath__24_0_I1589 (.Y(N3036), .A(N2629));
OAI21XL inst_cellmath__24_0_I1590 (.Y(N3376), .A0(N2669), .A1(N3522), .B0(N3036));
AOI21XL inst_cellmath__24_0_I1591 (.Y(N3176), .A0(N2787), .A1(N3306), .B0(N2423));
AOI21XL inst_cellmath__24_0_I1592 (.Y(N2972), .A0(N2571), .A1(N3325), .B0(N2219));
AOI21XL inst_cellmath__24_0_I1593 (.Y(N2761), .A0(N2360), .A1(N3643), .B0(N3623));
AOI21XL inst_cellmath__24_0_I1594 (.Y(N2550), .A0(N2161), .A1(N3121), .B0(N3422));
AOI21XL inst_cellmath__24_0_I1595 (.Y(N2336), .A0(N3564), .A1(N2383), .B0(N3225));
AOI21XL inst_cellmath__24_0_I1596 (.Y(N3746), .A0(N3367), .A1(N2914), .B0(N3025));
AOI21XL inst_cellmath__24_0_I1597 (.Y(N3542), .A0(N3166), .A1(N2707), .B0(N2811));
XNOR2X1 inst_cellmath__24_0_I1598 (.Y(inst_cellmath__24[19]), .A(N2459), .B(N3513));
XOR2XL inst_cellmath__24_0_I1599 (.Y(inst_cellmath__24[20]), .A(N2600), .B(N2606));
XNOR2X1 inst_cellmath__24_0_I1600 (.Y(inst_cellmath__24[21]), .A(N2495), .B(N3314));
XNOR2X1 inst_cellmath__24_0_I1601 (.Y(inst_cellmath__24[22]), .A(N3471), .B(N2396));
XOR2XL inst_cellmath__24_0_I1602 (.Y(inst_cellmath__24[23]), .A(N2285), .B(N3112));
XOR2XL inst_cellmath__24_0_I1603 (.Y(inst_cellmath__24[24]), .A(N3242), .B(N2193));
XNOR2X1 inst_cellmath__24_0_I1604 (.Y(inst_cellmath__24[25]), .A(N2798), .B(N2904));
XNOR2X1 inst_cellmath__24_0_I1605 (.Y(inst_cellmath__24[26]), .A(N2595), .B(N3596));
XOR2XL inst_cellmath__24_0_I1606 (.Y(inst_cellmath__24[27]), .A(N2584), .B(N2692));
XNOR2X1 inst_cellmath__24_0_I1607 (.Y(inst_cellmath__24[28]), .A(N3044), .B(N3395));
XOR2XL inst_cellmath__24_0_I1608 (.Y(inst_cellmath__24[29]), .A(N2367), .B(N2483));
XOR2XL inst_cellmath__24_0_I1609 (.Y(inst_cellmath__24[30]), .A(N2958), .B(N3197));
XNOR2X1 inst_cellmath__24_0_I1610 (.Y(inst_cellmath__24[31]), .A(N2879), .B(N2274));
XOR2XL inst_cellmath__24_0_I1611 (.Y(inst_cellmath__24[32]), .A(N3522), .B(N2995));
XNOR2X1 inst_cellmath__24_0_I1612 (.Y(inst_cellmath__24[33]), .A(N3376), .B(N3680));
XNOR2X1 inst_cellmath__24_0_I1613 (.Y(inst_cellmath__24[34]), .A(N3306), .B(N2787));
XOR2XL inst_cellmath__24_0_I1614 (.Y(inst_cellmath__24[35]), .A(N3176), .B(N3480));
XNOR2X1 inst_cellmath__24_0_I1615 (.Y(inst_cellmath__24[36]), .A(N3325), .B(N2571));
XOR2XL inst_cellmath__24_0_I1616 (.Y(inst_cellmath__24[37]), .A(N2972), .B(N3284));
XNOR2X1 inst_cellmath__24_0_I1617 (.Y(inst_cellmath__24[38]), .A(N3643), .B(N2360));
XOR2XL inst_cellmath__24_0_I1618 (.Y(inst_cellmath__24[39]), .A(N2761), .B(N3082));
XNOR2X1 inst_cellmath__24_0_I1619 (.Y(inst_cellmath__24[40]), .A(N3121), .B(N2161));
XOR2XL inst_cellmath__24_0_I1620 (.Y(inst_cellmath__24[41]), .A(N2550), .B(N2869));
XNOR2X1 inst_cellmath__24_0_I1621 (.Y(inst_cellmath__24[42]), .A(N2383), .B(N3564));
XOR2XL inst_cellmath__24_0_I1622 (.Y(inst_cellmath__24[43]), .A(N2336), .B(N2659));
XNOR2X1 inst_cellmath__24_0_I1623 (.Y(inst_cellmath__24[44]), .A(N2914), .B(N3367));
XOR2XL inst_cellmath__24_0_I1624 (.Y(inst_cellmath__24[45]), .A(N3746), .B(N2449));
XNOR2X1 inst_cellmath__24_0_I1625 (.Y(inst_cellmath__24[46]), .A(N2707), .B(N3166));
XNOR2X1 inst_cellmath__24_0_I1626 (.Y(inst_cellmath__24[47]), .A(N3542), .B(N2244));
BUFX2 inst_cellmath__25_0_I1627 (.Y(N5360), .A(inst_cellmath__24[47]));
AND2XL inst_cellmath__25_0_I1628 (.Y(inst_cellmath__25[0]), .A(N5360), .B(inst_cellmath__24[0]));
MX2XL inst_cellmath__25_0_I1629 (.Y(inst_cellmath__25[1]), .A(inst_cellmath__24[0]), .B(inst_cellmath__24[1]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1630 (.Y(inst_cellmath__25[2]), .A(inst_cellmath__24[1]), .B(inst_cellmath__24[2]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1631 (.Y(inst_cellmath__25[3]), .A(inst_cellmath__24[2]), .B(inst_cellmath__24[3]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1632 (.Y(inst_cellmath__25[4]), .A(inst_cellmath__24[3]), .B(inst_cellmath__24[4]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1633 (.Y(inst_cellmath__25[5]), .A(inst_cellmath__24[4]), .B(inst_cellmath__24[5]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1634 (.Y(inst_cellmath__25[6]), .A(inst_cellmath__24[5]), .B(inst_cellmath__24[6]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1635 (.Y(inst_cellmath__25[7]), .A(inst_cellmath__24[6]), .B(inst_cellmath__24[7]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1636 (.Y(inst_cellmath__25[8]), .A(inst_cellmath__24[7]), .B(inst_cellmath__24[8]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1637 (.Y(inst_cellmath__25[9]), .A(inst_cellmath__24[8]), .B(inst_cellmath__24[9]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1638 (.Y(inst_cellmath__25[10]), .A(inst_cellmath__24[9]), .B(inst_cellmath__24[10]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1639 (.Y(inst_cellmath__25[11]), .A(inst_cellmath__24[10]), .B(inst_cellmath__24[11]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1640 (.Y(inst_cellmath__25[12]), .A(inst_cellmath__24[11]), .B(inst_cellmath__24[12]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1641 (.Y(inst_cellmath__25[13]), .A(inst_cellmath__24[12]), .B(inst_cellmath__24[13]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1642 (.Y(inst_cellmath__25[14]), .A(inst_cellmath__24[13]), .B(inst_cellmath__24[14]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1643 (.Y(inst_cellmath__25[15]), .A(inst_cellmath__24[14]), .B(inst_cellmath__24[15]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1644 (.Y(inst_cellmath__25[16]), .A(inst_cellmath__24[15]), .B(inst_cellmath__24[16]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1645 (.Y(inst_cellmath__25[17]), .A(inst_cellmath__24[16]), .B(inst_cellmath__24[17]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1646 (.Y(inst_cellmath__25[18]), .A(inst_cellmath__24[17]), .B(inst_cellmath__24[18]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1647 (.Y(inst_cellmath__25[19]), .A(inst_cellmath__24[18]), .B(inst_cellmath__24[19]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1648 (.Y(inst_cellmath__25[20]), .A(inst_cellmath__24[19]), .B(inst_cellmath__24[20]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1649 (.Y(inst_cellmath__25[21]), .A(inst_cellmath__24[20]), .B(inst_cellmath__24[21]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1650 (.Y(inst_cellmath__25[22]), .A(inst_cellmath__24[21]), .B(inst_cellmath__24[22]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1651 (.Y(inst_cellmath__25[23]), .A(inst_cellmath__24[22]), .B(inst_cellmath__24[23]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1652 (.Y(inst_cellmath__25[24]), .A(inst_cellmath__24[23]), .B(inst_cellmath__24[24]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1653 (.Y(inst_cellmath__25[25]), .A(inst_cellmath__24[24]), .B(inst_cellmath__24[25]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1654 (.Y(inst_cellmath__25[26]), .A(inst_cellmath__24[25]), .B(inst_cellmath__24[26]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1655 (.Y(inst_cellmath__25[27]), .A(inst_cellmath__24[26]), .B(inst_cellmath__24[27]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1656 (.Y(inst_cellmath__25[28]), .A(inst_cellmath__24[27]), .B(inst_cellmath__24[28]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1657 (.Y(inst_cellmath__25[29]), .A(inst_cellmath__24[28]), .B(inst_cellmath__24[29]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1658 (.Y(inst_cellmath__25[30]), .A(inst_cellmath__24[29]), .B(inst_cellmath__24[30]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1659 (.Y(inst_cellmath__25[31]), .A(inst_cellmath__24[30]), .B(inst_cellmath__24[31]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1660 (.Y(inst_cellmath__25[32]), .A(inst_cellmath__24[31]), .B(inst_cellmath__24[32]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1661 (.Y(inst_cellmath__25[33]), .A(inst_cellmath__24[32]), .B(inst_cellmath__24[33]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1662 (.Y(inst_cellmath__25[34]), .A(inst_cellmath__24[33]), .B(inst_cellmath__24[34]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1663 (.Y(inst_cellmath__25[35]), .A(inst_cellmath__24[34]), .B(inst_cellmath__24[35]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1664 (.Y(inst_cellmath__25[36]), .A(inst_cellmath__24[35]), .B(inst_cellmath__24[36]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1665 (.Y(inst_cellmath__25[37]), .A(inst_cellmath__24[36]), .B(inst_cellmath__24[37]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1666 (.Y(inst_cellmath__25[38]), .A(inst_cellmath__24[37]), .B(inst_cellmath__24[38]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1667 (.Y(inst_cellmath__25[39]), .A(inst_cellmath__24[38]), .B(inst_cellmath__24[39]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1668 (.Y(inst_cellmath__25[40]), .A(inst_cellmath__24[39]), .B(inst_cellmath__24[40]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1669 (.Y(inst_cellmath__25[41]), .A(inst_cellmath__24[40]), .B(inst_cellmath__24[41]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1670 (.Y(inst_cellmath__25[42]), .A(inst_cellmath__24[41]), .B(inst_cellmath__24[42]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1671 (.Y(inst_cellmath__25[43]), .A(inst_cellmath__24[42]), .B(inst_cellmath__24[43]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1672 (.Y(inst_cellmath__25[44]), .A(inst_cellmath__24[43]), .B(inst_cellmath__24[44]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1673 (.Y(inst_cellmath__25[45]), .A(inst_cellmath__24[44]), .B(inst_cellmath__24[45]), .S0(N5360));
MX2XL inst_cellmath__25_0_I1674 (.Y(inst_cellmath__25[46]), .A(inst_cellmath__24[45]), .B(inst_cellmath__24[46]), .S0(N5360));
NOR2XL inst_cellmath__25_0_I1675 (.Y(inst_cellmath__25[47]), .A(N5360), .B(inst_cellmath__24[46]));
INVXL inst_cellmath__45_0_I1676 (.Y(inst_cellmath__45[0]), .A(inst_cellmath__25[24]));
NAND2XL inst_cellmath__45_0_I1677 (.Y(N5547), .A(inst_cellmath__25[26]), .B(inst_cellmath__25[25]));
NOR2XL inst_cellmath__45_0_I1678 (.Y(N5523), .A(N5547), .B(inst_cellmath__45[0]));
NAND2XL inst_cellmath__45_0_I1679 (.Y(N5552), .A(inst_cellmath__25[28]), .B(inst_cellmath__25[27]));
NAND4BXL inst_cellmath__45_0_I10379 (.Y(N5509), .AN(N5552), .B(inst_cellmath__25[30]), .C(N5523), .D(inst_cellmath__25[29]));
NAND2XL inst_cellmath__45_0_I1682 (.Y(N5511), .A(inst_cellmath__25[27]), .B(N5523));
NAND2BXL inst_cellmath__45_0_I1683 (.Y(N5482), .AN(N5552), .B(N5523));
NAND3BXL inst_cellmath__45_0_I1684 (.Y(N5542), .AN(N5552), .B(inst_cellmath__25[29]), .C(N5523));
NAND2XL inst_cellmath__45_0_I1686 (.Y(N5539), .A(inst_cellmath__25[32]), .B(inst_cellmath__25[31]));
NAND2XL inst_cellmath__45_0_I1687 (.Y(N5526), .A(inst_cellmath__25[34]), .B(inst_cellmath__25[33]));
NOR2XL inst_cellmath__45_0_I1688 (.Y(N5501), .A(N5526), .B(N5539));
NAND2XL inst_cellmath__45_0_I1689 (.Y(N5489), .A(inst_cellmath__25[36]), .B(inst_cellmath__25[35]));
NAND4BXL inst_cellmath__45_0_I10380 (.Y(N5496), .AN(N5489), .B(inst_cellmath__25[38]), .C(N5501), .D(inst_cellmath__25[37]));
NAND3BXL inst_cellmath__45_0_I1692 (.Y(N5554), .AN(N5489), .B(inst_cellmath__25[37]), .C(N5501));
NOR3BXL inst_cellmath__45_0_I1694 (.Y(N5499), .AN(inst_cellmath__25[33]), .B(N5539), .C(N5509));
NOR3BXL inst_cellmath__45_0_I1695 (.Y(N5495), .AN(N5501), .B(N5489), .C(N5509));
NOR2XL inst_cellmath__45_0_I1696 (.Y(N5528), .A(N5496), .B(N5509));
NAND2XL inst_cellmath__45_0_I1697 (.Y(N5557), .A(inst_cellmath__25[40]), .B(inst_cellmath__25[39]));
NAND2XL inst_cellmath__45_0_I1698 (.Y(N5544), .A(inst_cellmath__25[42]), .B(inst_cellmath__25[41]));
NOR2XL inst_cellmath__45_0_I1699 (.Y(N5520), .A(N5544), .B(N5557));
NAND2XL inst_cellmath__45_0_I1700 (.Y(N5507), .A(inst_cellmath__25[44]), .B(inst_cellmath__25[43]));
NAND2XL inst_cellmath__45_0_I1701 (.Y(N5506), .A(inst_cellmath__25[46]), .B(inst_cellmath__25[45]));
NOR2XL inst_cellmath__45_0_I1702 (.Y(N5473), .A(N5507), .B(N5506));
NAND2BXL inst_cellmath__45_0_I1705 (.Y(N5474), .AN(inst_cellmath__45[0]), .B(inst_cellmath__25[25]));
NAND2BXL inst_cellmath__45_0_I1706 (.Y(N5497), .AN(N5509), .B(inst_cellmath__25[31]));
OR2XL inst_cellmath__45_0_I1707 (.Y(N5521), .A(N5539), .B(N5509));
NAND2BXL inst_cellmath__45_0_I1708 (.Y(N5469), .AN(N5509), .B(N5501));
NAND3BXL inst_cellmath__45_0_I1709 (.Y(N5487), .AN(N5509), .B(inst_cellmath__25[35]), .C(N5501));
OR2XL inst_cellmath__45_0_I1710 (.Y(N5530), .A(N5554), .B(N5509));
NAND2XL inst_cellmath__45_0_I1711 (.Y(N5480), .A(inst_cellmath__25[39]), .B(N5528));
NAND2BXL inst_cellmath__45_0_I1712 (.Y(N5540), .AN(N5557), .B(N5528));
NAND3BXL inst_cellmath__45_0_I1713 (.Y(N5505), .AN(N5557), .B(inst_cellmath__25[41]), .C(N5528));
NAND2XL inst_cellmath__45_0_I1714 (.Y(N5477), .A(N5520), .B(N5528));
NAND3XL inst_cellmath__45_0_I1715 (.Y(N5536), .A(inst_cellmath__25[43]), .B(N5520), .C(N5528));
NAND3BXL inst_cellmath__45_0_I1716 (.Y(N5502), .AN(N5507), .B(N5520), .C(N5528));
NAND4BXL inst_cellmath__45_0_I1717 (.Y(N5472), .AN(N5507), .B(inst_cellmath__25[45]), .C(N5528), .D(N5520));
NAND3XL hyperpropagate_4_1_A_I3671 (.Y(N8442), .A(N5473), .B(N5528), .C(N5520));
NOR2XL hyperpropagate_4_1_A_I3672 (.Y(inst_cellmath__45[24]), .A(inst_cellmath__25[47]), .B(N8442));
XNOR2X1 inst_cellmath__45_0_I1720 (.Y(inst_cellmath__45[1]), .A(inst_cellmath__45[0]), .B(inst_cellmath__25[25]));
XNOR2X1 inst_cellmath__45_0_I1721 (.Y(inst_cellmath__45[2]), .A(N5474), .B(inst_cellmath__25[26]));
XOR2XL inst_cellmath__45_0_I1722 (.Y(inst_cellmath__45[3]), .A(N5523), .B(inst_cellmath__25[27]));
XNOR2X1 inst_cellmath__45_0_I1723 (.Y(inst_cellmath__45[4]), .A(N5511), .B(inst_cellmath__25[28]));
XNOR2X1 inst_cellmath__45_0_I1724 (.Y(inst_cellmath__45[5]), .A(N5482), .B(inst_cellmath__25[29]));
XNOR2X1 inst_cellmath__45_0_I1725 (.Y(inst_cellmath__45[6]), .A(N5542), .B(inst_cellmath__25[30]));
XNOR2X1 inst_cellmath__45_0_I1726 (.Y(inst_cellmath__45[7]), .A(N5509), .B(inst_cellmath__25[31]));
XNOR2X1 inst_cellmath__45_0_I1727 (.Y(inst_cellmath__45[8]), .A(N5497), .B(inst_cellmath__25[32]));
XNOR2X1 inst_cellmath__45_0_I1728 (.Y(inst_cellmath__45[9]), .A(N5521), .B(inst_cellmath__25[33]));
XOR2XL inst_cellmath__45_0_I1729 (.Y(inst_cellmath__45[10]), .A(N5499), .B(inst_cellmath__25[34]));
XNOR2X1 inst_cellmath__45_0_I1730 (.Y(inst_cellmath__45[11]), .A(N5469), .B(inst_cellmath__25[35]));
XNOR2X1 inst_cellmath__45_0_I1731 (.Y(inst_cellmath__45[12]), .A(N5487), .B(inst_cellmath__25[36]));
XOR2XL inst_cellmath__45_0_I1732 (.Y(inst_cellmath__45[13]), .A(N5495), .B(inst_cellmath__25[37]));
XNOR2X1 inst_cellmath__45_0_I1733 (.Y(inst_cellmath__45[14]), .A(N5530), .B(inst_cellmath__25[38]));
XOR2XL inst_cellmath__45_0_I1734 (.Y(inst_cellmath__45[15]), .A(N5528), .B(inst_cellmath__25[39]));
XNOR2X1 inst_cellmath__45_0_I1735 (.Y(inst_cellmath__45[16]), .A(N5480), .B(inst_cellmath__25[40]));
XNOR2X1 inst_cellmath__45_0_I1736 (.Y(inst_cellmath__45[17]), .A(N5540), .B(inst_cellmath__25[41]));
XNOR2X1 inst_cellmath__45_0_I1737 (.Y(inst_cellmath__45[18]), .A(N5505), .B(inst_cellmath__25[42]));
XNOR2X1 inst_cellmath__45_0_I1738 (.Y(inst_cellmath__45[19]), .A(N5477), .B(inst_cellmath__25[43]));
XNOR2X1 inst_cellmath__45_0_I1739 (.Y(inst_cellmath__45[20]), .A(N5536), .B(inst_cellmath__25[44]));
XNOR2X1 inst_cellmath__45_0_I1740 (.Y(inst_cellmath__45[21]), .A(N5502), .B(inst_cellmath__25[45]));
XNOR2X1 inst_cellmath__45_0_I1741 (.Y(inst_cellmath__45[22]), .A(N5472), .B(inst_cellmath__25[46]));
NOR3BXL cynw_cm_float_mul_ieee_I1743 (.Y(inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
INVXL inst_cellmath__44__31__I1744 (.Y(N5634), .A(inst_cellmath__23));
AND2XL inst_cellmath__44__31__I1745 (.Y(N446), .A(inst_cellmath__5), .B(N5634));
NOR3BXL cynw_cm_float_mul_ieee_I1746 (.Y(inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
AND2XL cynw_cm_float_mul_ieee_I1747 (.Y(N445), .A(inst_cellmath__6), .B(inst_cellmath__23));
NOR3BXL cynw_cm_float_mul_ieee_I1748 (.Y(inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR2XL inst_cellmath__34_0_I1754 (.Y(N5664), .A(inst_cellmath__25[3]), .B(inst_cellmath__25[22]));
NOR2XL inst_cellmath__34_0_I1755 (.Y(N5674), .A(inst_cellmath__25[20]), .B(inst_cellmath__25[18]));
OR4X1 inst_cellmath__34_0_I10381 (.Y(N5679), .A(inst_cellmath__25[13]), .B(inst_cellmath__25[17]), .C(inst_cellmath__25[15]), .D(inst_cellmath__25[19]));
OR4X1 inst_cellmath__34_0_I10382 (.Y(N5688), .A(inst_cellmath__25[5]), .B(inst_cellmath__25[9]), .C(inst_cellmath__25[7]), .D(inst_cellmath__25[11]));
OR4X1 inst_cellmath__34_0_I10383 (.Y(N5662), .A(inst_cellmath__25[10]), .B(inst_cellmath__25[14]), .C(inst_cellmath__25[12]), .D(inst_cellmath__25[16]));
OR4X1 inst_cellmath__34_0_I10384 (.Y(N5672), .A(inst_cellmath__25[2]), .B(inst_cellmath__25[6]), .C(inst_cellmath__25[4]), .D(inst_cellmath__25[8]));
NOR4X1 inst_cellmath__34_0_I1764 (.Y(N5692), .A(inst_cellmath__25[0]), .B(inst_cellmath__25[1]), .C(inst_cellmath__25[21]), .D(N5679));
NAND3XL inst_cellmath__34_0_I1766 (.Y(N5666), .A(N5664), .B(N5674), .C(N5692));
OR4X1 inst_cellmath__34_0_I10385 (.Y(inst_cellmath__34), .A(N5672), .B(N5662), .C(N5688), .D(N5666));
OR2XL cynw_cm_float_mul_ieee_I1769 (.Y(N443), .A(inst_cellmath__25[24]), .B(inst_cellmath__34));
NOR4BX1 cynw_cm_float_mul_ieee_I3655 (.Y(N444), .AN(N443), .B(rm[1]), .C(rm[0]), .D(rm[2]));
OR4X1 cynw_cm_float_mul_ieee_I1771 (.Y(N447), .A(inst_cellmath__8), .B(N445), .C(N446), .D(N444));
OAI21XL cynw_cm_float_mul_ieee_I3656 (.Y(N450), .A0(N445), .A1(N446), .B0(inst_cellmath__34));
OAI2BB1X1 cynw_cm_float_mul_ieee_I3657 (.Y(inst_cellmath__44), .A0N(inst_cellmath__25[23]), .A1N(N447), .B0(N450));
AOI21XL cynw_cm_float_mul_ieee_I3658 (.Y(inst_cellmath__38), .A0(inst_cellmath__45[24]), .A1(inst_cellmath__44), .B0(inst_cellmath__24[47]));
INVXL inst_cellmath__30_0_I1778 (.Y(N5761), .A(a_exp[7]));
XNOR2X1 inst_cellmath__30_0_I1779 (.Y(inst_cellmath__30[0]), .A(b_exp[0]), .B(a_exp[0]));
OR2XL inst_cellmath__30_0_I1780 (.Y(N5765), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 inst_cellmath__30_0_I1781 (.CO(N5758), .S(inst_cellmath__30[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(N5765));
ADDFX1 inst_cellmath__30_0_I1782 (.CO(N5777), .S(inst_cellmath__30[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(N5758));
ADDFX1 inst_cellmath__30_0_I1783 (.CO(N5789), .S(inst_cellmath__30[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(N5777));
ADDFX1 inst_cellmath__30_0_I1784 (.CO(N5771), .S(inst_cellmath__30[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(N5789));
ADDFX1 inst_cellmath__30_0_I1785 (.CO(N5786), .S(inst_cellmath__30[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(N5771));
ADDFX1 inst_cellmath__30_0_I1786 (.CO(N5766), .S(inst_cellmath__30[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(N5786));
ADDFX1 inst_cellmath__30_0_I1787 (.CO(N5781), .S(inst_cellmath__30[7]), .A(N5761), .B(b_exp[7]), .CI(N5766));
XNOR2X1 inst_cellmath__30_0_I1788 (.Y(inst_cellmath__30[8]), .A(a_exp[7]), .B(N5781));
NOR2XL inst_cellmath__30_0_I1789 (.Y(inst_cellmath__30[9]), .A(a_exp[7]), .B(N5781));
INVXL inst_cellmath__31_0_I1790 (.Y(inst_cellmath__31[0]), .A(inst_cellmath__30[0]));
NOR2BX1 inst_cellmath__31_0_I1791 (.Y(N5831), .AN(inst_cellmath__30[1]), .B(inst_cellmath__31[0]));
AND2XL inst_cellmath__31_0_I1792 (.Y(N5816), .A(inst_cellmath__30[2]), .B(N5831));
XNOR2X1 inst_cellmath__31_0_I1793 (.Y(inst_cellmath__31[1]), .A(inst_cellmath__31[0]), .B(inst_cellmath__30[1]));
XOR2XL inst_cellmath__31_0_I1794 (.Y(inst_cellmath__31[2]), .A(N5831), .B(inst_cellmath__30[2]));
AND2XL inst_cellmath__31_0_I1795 (.Y(N5835), .A(inst_cellmath__30[3]), .B(N5816));
AND3XL inst_cellmath__31_0_I1796 (.Y(N5834), .A(inst_cellmath__30[4]), .B(inst_cellmath__30[5]), .C(N5835));
AND3XL inst_cellmath__31_0_I1797 (.Y(N5825), .A(inst_cellmath__30[6]), .B(inst_cellmath__30[7]), .C(N5834));
NAND2XL inst_cellmath__31_0_I1798 (.Y(N5815), .A(inst_cellmath__30[4]), .B(N5835));
NAND2XL inst_cellmath__31_0_I1799 (.Y(N5833), .A(inst_cellmath__30[6]), .B(N5834));
NAND2XL inst_cellmath__31_0_I1800 (.Y(N5824), .A(inst_cellmath__30[8]), .B(N5825));
XOR2XL inst_cellmath__31_0_I1801 (.Y(inst_cellmath__31[3]), .A(N5816), .B(inst_cellmath__30[3]));
XOR2XL inst_cellmath__31_0_I1802 (.Y(inst_cellmath__31[4]), .A(N5835), .B(inst_cellmath__30[4]));
XNOR2X1 inst_cellmath__31_0_I1803 (.Y(inst_cellmath__31[5]), .A(N5815), .B(inst_cellmath__30[5]));
XOR2XL inst_cellmath__31_0_I1804 (.Y(inst_cellmath__31[6]), .A(N5834), .B(inst_cellmath__30[6]));
XNOR2X1 inst_cellmath__31_0_I1805 (.Y(inst_cellmath__31[7]), .A(N5833), .B(inst_cellmath__30[7]));
XOR2XL inst_cellmath__31_0_I1806 (.Y(inst_cellmath__31[8]), .A(N5825), .B(inst_cellmath__30[8]));
XNOR2X1 inst_cellmath__31_0_I1807 (.Y(inst_cellmath__31[9]), .A(N5824), .B(inst_cellmath__30[9]));
MX2XL inst_cellmath__48_0_I1808 (.Y(inst_cellmath__48[0]), .A(inst_cellmath__31[0]), .B(inst_cellmath__30[0]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1809 (.Y(inst_cellmath__48[1]), .A(inst_cellmath__31[1]), .B(inst_cellmath__30[1]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1810 (.Y(inst_cellmath__48[2]), .A(inst_cellmath__31[2]), .B(inst_cellmath__30[2]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1811 (.Y(inst_cellmath__48[3]), .A(inst_cellmath__31[3]), .B(inst_cellmath__30[3]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1812 (.Y(inst_cellmath__48[4]), .A(inst_cellmath__31[4]), .B(inst_cellmath__30[4]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1813 (.Y(inst_cellmath__48[5]), .A(inst_cellmath__31[5]), .B(inst_cellmath__30[5]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1814 (.Y(inst_cellmath__48[6]), .A(inst_cellmath__31[6]), .B(inst_cellmath__30[6]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1815 (.Y(inst_cellmath__48[7]), .A(inst_cellmath__31[7]), .B(inst_cellmath__30[7]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1816 (.Y(inst_cellmath__48[8]), .A(inst_cellmath__31[8]), .B(inst_cellmath__30[8]), .S0(inst_cellmath__38));
MX2XL inst_cellmath__48_0_I1817 (.Y(inst_cellmath__48[9]), .A(inst_cellmath__31[9]), .B(inst_cellmath__30[9]), .S0(inst_cellmath__38));
NAND2XL inst_cellmath__51__49__I1819 (.Y(N5906), .A(inst_cellmath__48[0]), .B(inst_cellmath__48[5]));
NAND2XL inst_cellmath__51__49__I1820 (.Y(N5909), .A(inst_cellmath__48[4]), .B(inst_cellmath__48[2]));
NAND2XL inst_cellmath__51__49__I1821 (.Y(N5897), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[3]));
NOR2XL inst_cellmath__51__49__I1823 (.Y(N5904), .A(N5909), .B(N5897));
NAND3XL hyperpropagate_4_1_A_I3673 (.Y(N8450), .A(inst_cellmath__48[1]), .B(inst_cellmath__48[6]), .C(N5904));
NOR2XL hyperpropagate_4_1_A_I3674 (.Y(N461), .A(N5906), .B(N8450));
NOR2XL andori2bb1_A_I3675 (.Y(N8456), .A(inst_cellmath__48[8]), .B(N461));
NOR2XL andori2bb1_A_I3676 (.Y(inst_cellmath__51), .A(N8456), .B(inst_cellmath__48[9]));
NAND2XL cynw_cm_float_mul_ieee_I1827 (.Y(inst_cellmath__28), .A(inst_cellmath__20), .B(inst_cellmath__13));
NAND2XL cynw_cm_float_mul_ieee_I1828 (.Y(inst_cellmath__27), .A(inst_cellmath__21), .B(inst_cellmath__14));
OR4X1 inst_cellmath__50__50__I10387 (.Y(N5949), .A(inst_cellmath__48[8]), .B(inst_cellmath__48[6]), .C(inst_cellmath__48[1]), .D(inst_cellmath__48[9]));
NOR4X1 inst_cellmath__50__50__I1832 (.Y(N5946), .A(inst_cellmath__48[0]), .B(inst_cellmath__48[2]), .C(inst_cellmath__48[4]), .D(inst_cellmath__48[5]));
NOR3XL inst_cellmath__50__50__I1833 (.Y(N5942), .A(inst_cellmath__48[7]), .B(inst_cellmath__48[3]), .C(N5949));
NOR4X1 inst_cellmath__49_1_I1835 (.Y(N5964), .A(inst_cellmath__28), .B(inst_cellmath__27), .C(inst_cellmath__26), .D(inst_cellmath__48[9]));
OAI2BB1X1 inst_cellmath__49_1_I3661 (.Y(N5957), .A0N(N5946), .A1N(N5942), .B0(N5964));
OR2XL inst_cellmath__49_1_I1837 (.Y(inst_cellmath__49), .A(N5957), .B(inst_cellmath__51));
OR2XL cynw_cm_float_mul_ieee_I1838 (.Y(N470), .A(inst_cellmath__27), .B(inst_cellmath__26));
OR2XL cynw_cm_float_mul_ieee_I1839 (.Y(N442), .A(inst_cellmath__30[8]), .B(inst_cellmath__30[7]));
NAND2BXL cynw_cm_float_mul_ieee_I1840 (.Y(inst_cellmath__32), .AN(inst_cellmath__30[9]), .B(N442));
NOR2XL cynw_cm_float_mul_ieee_I1841 (.Y(N469), .A(inst_cellmath__28), .B(inst_cellmath__32));
NAND2XL inst_cellmath__7_0_I1842 (.Y(N5986), .A(rm[0]), .B(rm[1]));
NOR2XL inst_cellmath__7_0_I1843 (.Y(inst_cellmath__7), .A(rm[2]), .B(N5986));
MXI2XL inst_cellmath__42_0_I1845 (.Y(N5994), .A(inst_cellmath__7), .B(N5634), .S0(inst_cellmath__6));
MX2XL inst_cellmath__42_0_I1846 (.Y(inst_cellmath__42), .A(N5994), .B(N5634), .S0(inst_cellmath__5));
AOI21XL inst_cellmath__52_0_I1848 (.Y(N6025), .A0(inst_cellmath__42), .A1(N469), .B0(N470));
OR2XL inst_cellmath__52_0_I1849 (.Y(N6008), .A(N469), .B(N470));
INVXL inst_cellmath__52_0_I1850 (.Y(N6004), .A(inst_cellmath__48[0]));
MXI2XL inst_cellmath__52_0_I1851 (.Y(x[23]), .A(N6004), .B(N6025), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1852 (.Y(x[24]), .A(inst_cellmath__48[1]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1853 (.Y(x[25]), .A(inst_cellmath__48[2]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1854 (.Y(x[26]), .A(inst_cellmath__48[3]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1855 (.Y(x[27]), .A(inst_cellmath__48[4]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1856 (.Y(x[28]), .A(inst_cellmath__48[5]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1857 (.Y(x[29]), .A(inst_cellmath__48[6]), .B(N6008), .S0(inst_cellmath__49));
MX2XL inst_cellmath__52_0_I1858 (.Y(x[30]), .A(inst_cellmath__48[7]), .B(N6008), .S0(inst_cellmath__49));
OR4X1 inst_cellmath__47_0_I1859 (.Y(N6044), .A(inst_cellmath__28), .B(inst_cellmath__27), .C(inst_cellmath__26), .D(inst_cellmath__42));
NOR2XL inst_cellmath__47_0_I1860 (.Y(inst_cellmath__47), .A(N6044), .B(inst_cellmath__32));
NOR2XL inst_cellmath__53_U_I1861 (.Y(N6055), .A(inst_cellmath__26), .B(inst_cellmath__47));
MXI2XL inst_cellmath__53_U_I1862 (.Y(N6053), .A(inst_cellmath__25[46]), .B(inst_cellmath__45[22]), .S0(inst_cellmath__44));
MXI2XL inst_cellmath__53_U_I1863 (.Y(x[22]), .A(N6053), .B(N6055), .S0(inst_cellmath__49));
INVXL inst_cellmath__53_M_I1864 (.Y(N6123), .A(inst_cellmath__49));
NOR2XL inst_cellmath__53_M_I1865 (.Y(N6106), .A(inst_cellmath__26), .B(N6123));
NAND3BXL inst_cellmath__53_M_I1866 (.Y(N6144), .AN(inst_cellmath__15), .B(inst_cellmath__22), .C(inst_cellmath__26));
NOR2XL inst_cellmath__53_M_I1867 (.Y(N6192), .A(N6144), .B(N6123));
NAND2XL inst_cellmath__53_M_I1868 (.Y(N6225), .A(inst_cellmath__15), .B(inst_cellmath__26));
NOR2XL inst_cellmath__53_M_I1869 (.Y(N6082), .A(N6225), .B(N6123));
NOR2BX1 inst_cellmath__53_M_I1870 (.Y(N6117), .AN(N6123), .B(inst_cellmath__44));
AND2XL inst_cellmath__53_M_I1871 (.Y(N6158), .A(inst_cellmath__44), .B(N6123));
AOI22XL inst_cellmath__53_M_I1872 (.Y(N6244), .A0(inst_cellmath__45[0]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[24]));
AOI22XL inst_cellmath__53_M_I1873 (.Y(N6138), .A0(inst_cellmath__45[1]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[25]));
AOI22XL inst_cellmath__53_M_I1874 (.Y(N6218), .A0(inst_cellmath__45[2]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[26]));
AOI22XL inst_cellmath__53_M_I1875 (.Y(N6112), .A0(inst_cellmath__45[3]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[27]));
AOI22XL inst_cellmath__53_M_I1876 (.Y(N6196), .A0(inst_cellmath__45[4]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[28]));
AOI22XL inst_cellmath__53_M_I1877 (.Y(N6087), .A0(inst_cellmath__45[5]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[29]));
AOI22XL inst_cellmath__53_M_I1878 (.Y(N6170), .A0(inst_cellmath__45[6]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[30]));
AOI22XL inst_cellmath__53_M_I1879 (.Y(N6063), .A0(inst_cellmath__45[7]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[31]));
AOI22XL inst_cellmath__53_M_I1880 (.Y(N6148), .A0(inst_cellmath__45[8]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[32]));
AOI22XL inst_cellmath__53_M_I1881 (.Y(N6230), .A0(inst_cellmath__45[9]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[33]));
AOI22XL inst_cellmath__53_M_I1882 (.Y(N6122), .A0(inst_cellmath__45[10]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[34]));
AOI22XL inst_cellmath__53_M_I1883 (.Y(N6207), .A0(inst_cellmath__45[11]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[35]));
AOI22XL inst_cellmath__53_M_I1884 (.Y(N6097), .A0(inst_cellmath__45[12]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[36]));
AOI22XL inst_cellmath__53_M_I1885 (.Y(N6181), .A0(inst_cellmath__45[13]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[37]));
AOI22XL inst_cellmath__53_M_I1886 (.Y(N6071), .A0(inst_cellmath__45[14]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[38]));
AOI22XL inst_cellmath__53_M_I1887 (.Y(N6157), .A0(inst_cellmath__45[15]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[39]));
AOI22XL inst_cellmath__53_M_I1888 (.Y(N6239), .A0(inst_cellmath__45[16]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[40]));
AOI22XL inst_cellmath__53_M_I1889 (.Y(N6132), .A0(inst_cellmath__45[17]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[41]));
AOI22XL inst_cellmath__53_M_I1890 (.Y(N6214), .A0(inst_cellmath__45[18]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[42]));
AOI22XL inst_cellmath__53_M_I1891 (.Y(N6107), .A0(inst_cellmath__45[19]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[43]));
AOI22XL inst_cellmath__53_M_I1892 (.Y(N6191), .A0(inst_cellmath__45[20]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[44]));
AOI22XL inst_cellmath__53_M_I1893 (.Y(N6081), .A0(inst_cellmath__45[21]), .A1(N6158), .B0(N6117), .B1(inst_cellmath__25[45]));
AOI22XL inst_cellmath__53_M_I1894 (.Y(N6114), .A0(b_man[0]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1895 (.Y(N6089), .A0(b_man[1]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1896 (.Y(N6064), .A0(b_man[2]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1897 (.Y(N6232), .A0(b_man[3]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1898 (.Y(N6209), .A0(b_man[4]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1899 (.Y(N6183), .A0(b_man[5]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1900 (.Y(N6160), .A0(b_man[6]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1901 (.Y(N6134), .A0(b_man[7]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1902 (.Y(N6108), .A0(b_man[8]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1903 (.Y(N6083), .A0(b_man[9]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1904 (.Y(N6060), .A0(b_man[10]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1905 (.Y(N6226), .A0(b_man[11]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1906 (.Y(N6203), .A0(b_man[12]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1907 (.Y(N6177), .A0(b_man[13]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1908 (.Y(N6154), .A0(b_man[14]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1909 (.Y(N6129), .A0(b_man[15]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1910 (.Y(N6103), .A0(b_man[16]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1911 (.Y(N6078), .A0(b_man[17]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1912 (.Y(N6247), .A0(b_man[18]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1913 (.Y(N6221), .A0(b_man[19]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1914 (.Y(N6199), .A0(b_man[20]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
AOI22XL inst_cellmath__53_M_I1915 (.Y(N6173), .A0(b_man[21]), .A1(N6192), .B0(N6106), .B1(inst_cellmath__47));
NAND2XL inst_cellmath__53_M_I1916 (.Y(N6150), .A(N6082), .B(a_man[0]));
NAND2XL inst_cellmath__53_M_I1917 (.Y(N6234), .A(N6082), .B(a_man[1]));
NAND2XL inst_cellmath__53_M_I1918 (.Y(N6126), .A(N6082), .B(a_man[2]));
NAND2XL inst_cellmath__53_M_I1919 (.Y(N6210), .A(N6082), .B(a_man[3]));
NAND2XL inst_cellmath__53_M_I1920 (.Y(N6100), .A(N6082), .B(a_man[4]));
NAND2XL inst_cellmath__53_M_I1921 (.Y(N6185), .A(N6082), .B(a_man[5]));
NAND2XL inst_cellmath__53_M_I1922 (.Y(N6073), .A(N6082), .B(a_man[6]));
NAND2XL inst_cellmath__53_M_I1923 (.Y(N6162), .A(N6082), .B(a_man[7]));
NAND2XL inst_cellmath__53_M_I1924 (.Y(N6242), .A(N6082), .B(a_man[8]));
NAND2XL inst_cellmath__53_M_I1925 (.Y(N6135), .A(N6082), .B(a_man[9]));
NAND2XL inst_cellmath__53_M_I1926 (.Y(N6216), .A(N6082), .B(a_man[10]));
NAND2XL inst_cellmath__53_M_I1927 (.Y(N6110), .A(N6082), .B(a_man[11]));
NAND2XL inst_cellmath__53_M_I1928 (.Y(N6193), .A(N6082), .B(a_man[12]));
NAND2XL inst_cellmath__53_M_I1929 (.Y(N6085), .A(N6082), .B(a_man[13]));
NAND2XL inst_cellmath__53_M_I1930 (.Y(N6168), .A(N6082), .B(a_man[14]));
NAND2XL inst_cellmath__53_M_I1931 (.Y(N6061), .A(N6082), .B(a_man[15]));
NAND2XL inst_cellmath__53_M_I1932 (.Y(N6146), .A(N6082), .B(a_man[16]));
NAND2XL inst_cellmath__53_M_I1933 (.Y(N6228), .A(N6082), .B(a_man[17]));
NAND2XL inst_cellmath__53_M_I1934 (.Y(N6120), .A(N6082), .B(a_man[18]));
NAND2XL inst_cellmath__53_M_I1935 (.Y(N6205), .A(N6082), .B(a_man[19]));
NAND2XL inst_cellmath__53_M_I1936 (.Y(N6095), .A(N6082), .B(a_man[20]));
NAND2XL inst_cellmath__53_M_I1937 (.Y(N6178), .A(N6082), .B(a_man[21]));
NAND3XL inst_cellmath__53_M_I1938 (.Y(x[0]), .A(N6150), .B(N6244), .C(N6114));
NAND3XL inst_cellmath__53_M_I1939 (.Y(x[1]), .A(N6234), .B(N6138), .C(N6089));
NAND3XL inst_cellmath__53_M_I1940 (.Y(x[2]), .A(N6126), .B(N6218), .C(N6064));
NAND3XL inst_cellmath__53_M_I1941 (.Y(x[3]), .A(N6210), .B(N6112), .C(N6232));
NAND3XL inst_cellmath__53_M_I1942 (.Y(x[4]), .A(N6100), .B(N6196), .C(N6209));
NAND3XL inst_cellmath__53_M_I1943 (.Y(x[5]), .A(N6185), .B(N6087), .C(N6183));
NAND3XL inst_cellmath__53_M_I1944 (.Y(x[6]), .A(N6073), .B(N6170), .C(N6160));
NAND3XL inst_cellmath__53_M_I1945 (.Y(x[7]), .A(N6162), .B(N6063), .C(N6134));
NAND3XL inst_cellmath__53_M_I1946 (.Y(x[8]), .A(N6242), .B(N6148), .C(N6108));
NAND3XL inst_cellmath__53_M_I1947 (.Y(x[9]), .A(N6135), .B(N6230), .C(N6083));
NAND3XL inst_cellmath__53_M_I1948 (.Y(x[10]), .A(N6216), .B(N6122), .C(N6060));
NAND3XL inst_cellmath__53_M_I1949 (.Y(x[11]), .A(N6110), .B(N6207), .C(N6226));
NAND3XL inst_cellmath__53_M_I1950 (.Y(x[12]), .A(N6193), .B(N6097), .C(N6203));
NAND3XL inst_cellmath__53_M_I1951 (.Y(x[13]), .A(N6085), .B(N6181), .C(N6177));
NAND3XL inst_cellmath__53_M_I1952 (.Y(x[14]), .A(N6168), .B(N6071), .C(N6154));
NAND3XL inst_cellmath__53_M_I1953 (.Y(x[15]), .A(N6061), .B(N6157), .C(N6129));
NAND3XL inst_cellmath__53_M_I1954 (.Y(x[16]), .A(N6146), .B(N6239), .C(N6103));
NAND3XL inst_cellmath__53_M_I1955 (.Y(x[17]), .A(N6228), .B(N6132), .C(N6078));
NAND3XL inst_cellmath__53_M_I1956 (.Y(x[18]), .A(N6120), .B(N6214), .C(N6247));
NAND3XL inst_cellmath__53_M_I1957 (.Y(x[19]), .A(N6205), .B(N6107), .C(N6221));
NAND3XL inst_cellmath__53_M_I1958 (.Y(x[20]), .A(N6095), .B(N6191), .C(N6199));
NAND3XL inst_cellmath__53_M_I1959 (.Y(x[21]), .A(N6178), .B(N6081), .C(N6173));
assign inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  urf3SgnYrR0= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



