/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:10:30 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_0_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__9,
	inst_cellmath__17;
wire [8:0] inst_cellmath__19;
wire [7:0] inst_cellmath__20;
wire [8:0] inst_cellmath__22;
wire  inst_cellmath__28,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__33,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42;
wire [15:0] inst_cellmath__48;
wire [18:0] inst_cellmath__51;
wire [24:0] inst_cellmath__60;
wire [39:0] inst_cellmath__62__W0, inst_cellmath__62__W1,
	inst_cellmath__63__W0, inst_cellmath__63__W1;
wire [39:0] inst_cellmath__64;
wire  inst_cellmath__67;
wire N446,N447,N448,N449,N450,N451,N452 
	,N453,N454,N455,N456,N457,N458,N477,N478 
	,N479,N480,N481,N482,N483,N484,N485,N486 
	,N487,N488,N489,N490,N491,N492,N493,N494 
	,N495,N496,N497,N498,N499,N500,N501;
cynw_cm_float_rcp_inst_cellmath__9_0_bdw1471647203_bdw cynw_cm_float_rcp_I0 (.inst_cellmath__9_0_out0(inst_cellmath__9), .inst_cellmath__9_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_rcp_inst_cellmath__15__5__bdw1471647203_bdw cynw_cm_float_rcp_I1 (.inst_cellmath__15__5__out0(inst_cellmath__19[0]), .inst_cellmath__15__5__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_rcp_inst_cellmath__29_0_bdw1471647203_bdw cynw_cm_float_rcp_I2 (.inst_cellmath__29_0_out0(inst_cellmath__29), .inst_cellmath__29_0_in0(inst_cellmath__9), .inst_cellmath__29_0_in1(inst_cellmath__19[0]));
cynw_cm_float_rcp_inst_cellmath__37_0_bdw1471647203_bdw cynw_cm_float_rcp_I3 (.inst_cellmath__37_0_out0(x[31]), .inst_cellmath__37_0_in0(inst_cellmath__29), .inst_cellmath__37_0_in1(a_sign));
cynw_cm_float_rcp_inst_cellmath__28_0_bdw1471647203_bdw cynw_cm_float_rcp_I4 (.inst_cellmath__28_0_out0(inst_cellmath__28), .inst_cellmath__28_0_in0(inst_cellmath__9), .inst_cellmath__28_0_in1(inst_cellmath__19[0]));
INVXL cynw_cm_float_rcp_I5 (.Y(inst_cellmath__20[0]), .A(a_exp[0]));
INVXL cynw_cm_float_rcp_I6 (.Y(inst_cellmath__20[1]), .A(a_exp[1]));
INVXL cynw_cm_float_rcp_I7 (.Y(inst_cellmath__20[2]), .A(a_exp[2]));
INVXL cynw_cm_float_rcp_I8 (.Y(inst_cellmath__20[3]), .A(a_exp[3]));
INVXL cynw_cm_float_rcp_I9 (.Y(inst_cellmath__20[4]), .A(a_exp[4]));
INVXL cynw_cm_float_rcp_I10 (.Y(inst_cellmath__20[5]), .A(a_exp[5]));
INVXL cynw_cm_float_rcp_I11 (.Y(inst_cellmath__20[6]), .A(a_exp[6]));
INVXL cynw_cm_float_rcp_I12 (.Y(inst_cellmath__20[7]), .A(a_exp[7]));
cynw_cm_float_rcp_inst_cellmath__22_0_bdw1471647203_bdw cynw_cm_float_rcp_I13 (.inst_cellmath__22_0_out0({inst_cellmath__22[8], inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}), .inst_cellmath__22_0_in0({inst_cellmath__20[7], inst_cellmath__20[6], inst_cellmath__20[5], inst_cellmath__20[4], inst_cellmath__20[3], inst_cellmath__20[2], inst_cellmath__20[1], inst_cellmath__20[0]}), .inst_cellmath__22_0_in1(inst_cellmath__19[0]));
cynw_cm_float_rcp_inst_cellmath__17__6__bdw1471647203_bdw cynw_cm_float_rcp_I14 (.inst_cellmath__17__6__out0({N446}), .inst_cellmath__17__6__in0({inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}));
cynw_cm_float_rcp_inst_cellmath__17_0_bdw1471647203_bdw cynw_cm_float_rcp_I15 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({inst_cellmath__22[8]}), .inst_cellmath__17_0_in1({N446}));
cynw_cm_float_rcp_inst_cellmath__30_0_bdw1471647203_bdw cynw_cm_float_rcp_I16 (.inst_cellmath__30_0_out0(inst_cellmath__30), .inst_cellmath__30_0_in0(inst_cellmath__9), .inst_cellmath__30_0_in1(inst_cellmath__17));
cynw_cm_float_rcp_inst_cellmath__33__7__bdw1471647203_bdw cynw_cm_float_rcp_I17 (.inst_cellmath__33__7__out0({N447}), .inst_cellmath__33__7__in0(inst_cellmath__30), .inst_cellmath__33__7__in1(inst_cellmath__28));
cynw_cm_float_rcp_inst_cellmath__33_0_bdw1471647203_bdw cynw_cm_float_rcp_I18 (.inst_cellmath__33_0_out0(inst_cellmath__33), .inst_cellmath__33_0_in0({N447}), .inst_cellmath__33_0_in1(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__34_0_bdw1471647203_bdw cynw_cm_float_rcp_I19 (.inst_cellmath__34_0_out0(inst_cellmath__34), .inst_cellmath__34_0_in0(inst_cellmath__29), .inst_cellmath__34_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_rcp_inst_cellmath__42__9__bdw1471647203_bdw cynw_cm_float_rcp_I20 (.inst_cellmath__42__9__out0(inst_cellmath__42), .inst_cellmath__42__9__in0(inst_cellmath__34), .inst_cellmath__42__9__in1(inst_cellmath__33), .inst_cellmath__42__9__in2(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__38_0_bdw1471647203_bdw cynw_cm_float_rcp_I21 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__34), .inst_cellmath__38_0_in1(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__43_0_bdw1471647203_bdw cynw_cm_float_rcp_I22 (.inst_cellmath__43_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__43_0_in0(inst_cellmath__42), .inst_cellmath__43_0_in1(inst_cellmath__38), .inst_cellmath__43_0_in2({inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}));
cynw_cm_float_rcp_inst_cellmath__67__11__bdw1471647203_bdw cynw_cm_float_rcp_I23 (.inst_cellmath__67__11__out0({N448}), .inst_cellmath__67__11__in0(inst_cellmath__34), .inst_cellmath__67__11__in1(inst_cellmath__33), .inst_cellmath__67__11__in2(inst_cellmath__29), .inst_cellmath__67__11__in3(inst_cellmath__19[0]));
INVXL cynw_cm_float_rcp_I24 (.Y(inst_cellmath__67), .A(N448));
INVX1 cynw_cm_float_rcp_I25 (.Y(inst_cellmath__48[15]), .A(a_man[15]));
cynw_cm_float_rcp_inst_cellmath__60_0_bdw1471647203_bdw cynw_cm_float_rcp_I26 (.inst_cellmath__60_0_out0({inst_cellmath__60[24], inst_cellmath__60[23], inst_cellmath__60[22], inst_cellmath__60[21], inst_cellmath__60[20], inst_cellmath__60[19], inst_cellmath__60[18], inst_cellmath__60[17], inst_cellmath__60[16], inst_cellmath__60[15], inst_cellmath__60[14], inst_cellmath__60[13], inst_cellmath__60[12], inst_cellmath__60[11], inst_cellmath__60[10], inst_cellmath__60[9], inst_cellmath__60[8], inst_cellmath__60[7], inst_cellmath__60[6], inst_cellmath__60[5], inst_cellmath__60[4], inst_cellmath__60[3], inst_cellmath__60[2], inst_cellmath__60[1], inst_cellmath__60[0]}), .inst_cellmath__60_0_in0(inst_cellmath__48[15]), .inst_cellmath__60_0_in1({a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3]}));
cynw_cm_float_rcp_inst_noninc_a_cellmath__55_2WWMM_bdw1471647203_bdw cynw_cm_float_rcp_I27 (.inst_noninc_a_cellmath__55_2WWMM_out0({N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, inst_cellmath__51[17], inst_cellmath__51[16], inst_cellmath__51[15], inst_cellmath__51[14], inst_cellmath__51[13], inst_cellmath__51[12], inst_cellmath__51[11], inst_cellmath__51[10], inst_cellmath__51[9], inst_cellmath__51[8], inst_cellmath__51[7], inst_cellmath__51[6], inst_cellmath__51[5], inst_cellmath__51[4], inst_cellmath__51[3], inst_cellmath__51[2], inst_cellmath__51[1], inst_cellmath__51[0], N458, N457, N456, N455, N454, N453, N452, N451, N450, N449}), .inst_noninc_a_cellmath__55_2WWMM_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16]}));
cynw_cm_float_rcp_inst_cellmath__62_0_bdw1471647203_bdw cynw_cm_float_rcp_I28 (.inst_cellmath__62_0_out0({inst_cellmath__62__W1[39], inst_cellmath__62__W1[38], inst_cellmath__62__W1[37], inst_cellmath__62__W1[36], inst_cellmath__62__W1[35], inst_cellmath__62__W1[34], inst_cellmath__62__W1[33], inst_cellmath__62__W1[32], inst_cellmath__62__W1[31], inst_cellmath__62__W1[30], inst_cellmath__62__W1[29], inst_cellmath__62__W1[28], inst_cellmath__62__W1[27], inst_cellmath__62__W1[26], inst_cellmath__62__W1[25], inst_cellmath__62__W1[24], inst_cellmath__62__W1[23], inst_cellmath__62__W1[22], inst_cellmath__62__W1[21], inst_cellmath__62__W1[20], inst_cellmath__62__W1[19], inst_cellmath__62__W1[18], inst_cellmath__62__W1[17], inst_cellmath__62__W1[16], inst_cellmath__62__W1[15], inst_cellmath__62__W1[14], inst_cellmath__62__W1[13], inst_cellmath__62__W1[12], inst_cellmath__62__W1[11], inst_cellmath__62__W1[10], inst_cellmath__62__W1[9], inst_cellmath__62__W1[8], inst_cellmath__62__W1[7], inst_cellmath__62__W1[6], inst_cellmath__62__W1[5], inst_cellmath__62__W1[4], inst_cellmath__62__W1[3], inst_cellmath__62__W1[2], inst_cellmath__62__W1[1], inst_cellmath__62__W1[0]}), .inst_cellmath__62_0_out1({inst_cellmath__62__W0[39], inst_cellmath__62__W0[38], inst_cellmath__62__W0[37], inst_cellmath__62__W0[36], inst_cellmath__62__W0[35], inst_cellmath__62__W0[34], inst_cellmath__62__W0[33], inst_cellmath__62__W0[32], inst_cellmath__62__W0[31], inst_cellmath__62__W0[30], inst_cellmath__62__W0[29], inst_cellmath__62__W0[28], inst_cellmath__62__W0[27], inst_cellmath__62__W0[26], inst_cellmath__62__W0[25], inst_cellmath__62__W0[24], inst_cellmath__62__W0[23], inst_cellmath__62__W0[22], inst_cellmath__62__W0[21], inst_cellmath__62__W0[20], inst_cellmath__62__W0[19], inst_cellmath__62__W0[18], inst_cellmath__62__W0[17], inst_cellmath__62__W0[16], inst_cellmath__62__W0[15], inst_cellmath__62__W0[14], inst_cellmath__62__W0[13], inst_cellmath__62__W0[12], inst_cellmath__62__W0[11], inst_cellmath__62__W0[10], inst_cellmath__62__W0[9], inst_cellmath__62__W0[8], inst_cellmath__62__W0[7], inst_cellmath__62__W0[6], inst_cellmath__62__W0[5], inst_cellmath__62__W0[4], inst_cellmath__62__W0[3], inst_cellmath__62__W0[2], inst_cellmath__62__W0[1], inst_cellmath__62__W0[0]}), .inst_cellmath__62_0_in0({N458, N457, N456, N455, N454, N453, N452, N451, N450, N449}), .inst_cellmath__62_0_in1({inst_cellmath__60[24], inst_cellmath__60[23], inst_cellmath__60[22], inst_cellmath__60[21], inst_cellmath__60[20], inst_cellmath__60[19], inst_cellmath__60[18], inst_cellmath__60[17], inst_cellmath__60[16], inst_cellmath__60[15], inst_cellmath__60[14], inst_cellmath__60[13]}));
cynw_cm_float_rcp_inst_cellmath__63_0_bdw1471647203_bdw cynw_cm_float_rcp_I29 (.inst_cellmath__63_0_out0({inst_cellmath__63__W1[39], inst_cellmath__63__W1[38], inst_cellmath__63__W1[37], inst_cellmath__63__W1[36], inst_cellmath__63__W1[35], inst_cellmath__63__W1[34], inst_cellmath__63__W1[33], inst_cellmath__63__W1[32], inst_cellmath__63__W1[31], inst_cellmath__63__W1[30], inst_cellmath__63__W1[29], inst_cellmath__63__W1[28], inst_cellmath__63__W1[27], inst_cellmath__63__W1[26], inst_cellmath__63__W1[25], inst_cellmath__63__W1[24], inst_cellmath__63__W1[23], inst_cellmath__63__W1[22], inst_cellmath__63__W1[21], inst_cellmath__63__W1[20], inst_cellmath__63__W1[19], inst_cellmath__63__W1[18], inst_cellmath__63__W1[17], inst_cellmath__63__W1[16], inst_cellmath__63__W1[15], inst_cellmath__63__W1[14], inst_cellmath__63__W1[13], inst_cellmath__63__W1[12], inst_cellmath__63__W1[11], inst_cellmath__63__W1[10], inst_cellmath__63__W1[9], inst_cellmath__63__W1[8], inst_cellmath__63__W1[7], inst_cellmath__63__W1[6], inst_cellmath__63__W1[5], inst_cellmath__63__W1[4], inst_cellmath__63__W1[3], inst_cellmath__63__W1[2], inst_cellmath__63__W1[1], inst_cellmath__63__W1[0]}), .inst_cellmath__63_0_out1({inst_cellmath__63__W0[39], inst_cellmath__63__W0[38], inst_cellmath__63__W0[37], inst_cellmath__63__W0[36], inst_cellmath__63__W0[35], inst_cellmath__63__W0[34], inst_cellmath__63__W0[33], inst_cellmath__63__W0[32], inst_cellmath__63__W0[31], inst_cellmath__63__W0[30], inst_cellmath__63__W0[29], inst_cellmath__63__W0[28], inst_cellmath__63__W0[27], inst_cellmath__63__W0[26], inst_cellmath__63__W0[25], inst_cellmath__63__W0[24], inst_cellmath__63__W0[23], inst_cellmath__63__W0[22], inst_cellmath__63__W0[21], inst_cellmath__63__W0[20], inst_cellmath__63__W0[19], inst_cellmath__63__W0[18], inst_cellmath__63__W0[17], inst_cellmath__63__W0[16], inst_cellmath__63__W0[15], inst_cellmath__63__W0[14], inst_cellmath__63__W0[13], inst_cellmath__63__W0[12], inst_cellmath__63__W0[11], inst_cellmath__63__W0[10], inst_cellmath__63__W0[9], inst_cellmath__63__W0[8], inst_cellmath__63__W0[7], inst_cellmath__63__W0[6], inst_cellmath__63__W0[5], inst_cellmath__63__W0[4], inst_cellmath__63__W0[3], inst_cellmath__63__W0[2], inst_cellmath__63__W0[1], inst_cellmath__63__W0[0]}), .inst_cellmath__63_0_in0({inst_cellmath__51[17], inst_cellmath__51[16], inst_cellmath__51[15], inst_cellmath__51[14], inst_cellmath__51[13], inst_cellmath__51[12], inst_cellmath__51[11], inst_cellmath__51[10], inst_cellmath__51[9], inst_cellmath__51[8], inst_cellmath__51[7], inst_cellmath__51[6], inst_cellmath__51[5], inst_cellmath__51[4], inst_cellmath__51[3], inst_cellmath__51[2], inst_cellmath__51[1], inst_cellmath__51[0]}), .inst_cellmath__63_0_in1(inst_cellmath__48[15]), .inst_cellmath__63_0_in2({a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_rcp_inst_cellmath__64_0_bdw1471647203_bdw cynw_cm_float_rcp_I30 (.inst_cellmath__64_0_out0({inst_cellmath__64[39], inst_cellmath__64[38], inst_cellmath__64[37], inst_cellmath__64[36], inst_cellmath__64[35], inst_cellmath__64[34], inst_cellmath__64[33], inst_cellmath__64[32], inst_cellmath__64[31], inst_cellmath__64[30], inst_cellmath__64[29], inst_cellmath__64[28], inst_cellmath__64[27], inst_cellmath__64[26], inst_cellmath__64[25], inst_cellmath__64[24], inst_cellmath__64[23], inst_cellmath__64[22], inst_cellmath__64[21], inst_cellmath__64[20], inst_cellmath__64[19], inst_cellmath__64[18], inst_cellmath__64[17], inst_cellmath__64[16], inst_cellmath__64[15], inst_cellmath__64[14], inst_cellmath__64[13], inst_cellmath__64[12], inst_cellmath__64[11], inst_cellmath__64[10], inst_cellmath__64[9], inst_cellmath__64[8], inst_cellmath__64[7], inst_cellmath__64[6], inst_cellmath__64[5], inst_cellmath__64[4], inst_cellmath__64[3], inst_cellmath__64[2], inst_cellmath__64[1], inst_cellmath__64[0]}), .inst_cellmath__64_0_in0({N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477}), .inst_cellmath__64_0_in1({inst_cellmath__63__W1[39], inst_cellmath__63__W1[38], inst_cellmath__63__W1[37], inst_cellmath__63__W1[36], inst_cellmath__63__W1[35], inst_cellmath__63__W1[34], inst_cellmath__63__W1[33], inst_cellmath__63__W1[32], inst_cellmath__63__W1[31], inst_cellmath__63__W1[30], inst_cellmath__63__W1[29], inst_cellmath__63__W1[28], inst_cellmath__63__W1[27], inst_cellmath__63__W1[26], inst_cellmath__63__W1[25], inst_cellmath__63__W1[24], inst_cellmath__63__W1[23], inst_cellmath__63__W1[22], inst_cellmath__63__W1[21], inst_cellmath__63__W1[20], inst_cellmath__63__W1[19], inst_cellmath__63__W1[18], inst_cellmath__63__W1[17], inst_cellmath__63__W1[16], inst_cellmath__63__W1[15], inst_cellmath__63__W1[14], inst_cellmath__63__W1[13], inst_cellmath__63__W1[12], inst_cellmath__63__W1[11], inst_cellmath__63__W1[10], inst_cellmath__63__W1[9], inst_cellmath__63__W1[8], inst_cellmath__63__W1[7], inst_cellmath__63__W1[6], inst_cellmath__63__W1[5], inst_cellmath__63__W1[4], inst_cellmath__63__W1[3], inst_cellmath__63__W1[2], inst_cellmath__63__W1[1], inst_cellmath__63__W1[0]}), .inst_cellmath__64_0_in2({inst_cellmath__63__W0[39], inst_cellmath__63__W0[38], inst_cellmath__63__W0[37], inst_cellmath__63__W0[36], inst_cellmath__63__W0[35], inst_cellmath__63__W0[34], inst_cellmath__63__W0[33], inst_cellmath__63__W0[32], inst_cellmath__63__W0[31], inst_cellmath__63__W0[30], inst_cellmath__63__W0[29], inst_cellmath__63__W0[28], inst_cellmath__63__W0[27], inst_cellmath__63__W0[26], inst_cellmath__63__W0[25], inst_cellmath__63__W0[24], inst_cellmath__63__W0[23], inst_cellmath__63__W0[22], inst_cellmath__63__W0[21], inst_cellmath__63__W0[20], inst_cellmath__63__W0[19], inst_cellmath__63__W0[18], inst_cellmath__63__W0[17], inst_cellmath__63__W0[16], inst_cellmath__63__W0[15], inst_cellmath__63__W0[14], inst_cellmath__63__W0[13], inst_cellmath__63__W0[12], inst_cellmath__63__W0[11], inst_cellmath__63__W0[10], inst_cellmath__63__W0[9], inst_cellmath__63__W0[8], inst_cellmath__63__W0[7], inst_cellmath__63__W0[6], inst_cellmath__63__W0[5], inst_cellmath__63__W0[4], inst_cellmath__63__W0[3], inst_cellmath__63__W0[2], inst_cellmath__63__W0[1], inst_cellmath__63__W0[0]}), .inst_cellmath__64_0_in3({inst_cellmath__62__W1[39], inst_cellmath__62__W1[38], inst_cellmath__62__W1[37], inst_cellmath__62__W1[36], inst_cellmath__62__W1[35], inst_cellmath__62__W1[34], inst_cellmath__62__W1[33], inst_cellmath__62__W1[32], inst_cellmath__62__W1[31], inst_cellmath__62__W1[30], inst_cellmath__62__W1[29], inst_cellmath__62__W1[28], inst_cellmath__62__W1[27], inst_cellmath__62__W1[26], inst_cellmath__62__W1[25], inst_cellmath__62__W1[24], inst_cellmath__62__W1[23], inst_cellmath__62__W1[22], inst_cellmath__62__W1[21], inst_cellmath__62__W1[20], inst_cellmath__62__W1[19], inst_cellmath__62__W1[18], inst_cellmath__62__W1[17], inst_cellmath__62__W1[16], inst_cellmath__62__W1[15], inst_cellmath__62__W1[14], inst_cellmath__62__W1[13], inst_cellmath__62__W1[12], inst_cellmath__62__W1[11], inst_cellmath__62__W1[10], inst_cellmath__62__W1[9], inst_cellmath__62__W1[8], inst_cellmath__62__W1[7], inst_cellmath__62__W1[6], inst_cellmath__62__W1[5], inst_cellmath__62__W1[4], inst_cellmath__62__W1[3], inst_cellmath__62__W1[2], inst_cellmath__62__W1[1], inst_cellmath__62__W1[0]}), .inst_cellmath__64_0_in4({inst_cellmath__62__W0[39], inst_cellmath__62__W0[38], inst_cellmath__62__W0[37], inst_cellmath__62__W0[36], inst_cellmath__62__W0[35], inst_cellmath__62__W0[34], inst_cellmath__62__W0[33], inst_cellmath__62__W0[32], inst_cellmath__62__W0[31], inst_cellmath__62__W0[30], inst_cellmath__62__W0[29], inst_cellmath__62__W0[28], inst_cellmath__62__W0[27], inst_cellmath__62__W0[26], inst_cellmath__62__W0[25], inst_cellmath__62__W0[24], inst_cellmath__62__W0[23], inst_cellmath__62__W0[22], inst_cellmath__62__W0[21], inst_cellmath__62__W0[20], inst_cellmath__62__W0[19], inst_cellmath__62__W0[18], inst_cellmath__62__W0[17], inst_cellmath__62__W0[16], inst_cellmath__62__W0[15], inst_cellmath__62__W0[14], inst_cellmath__62__W0[13], inst_cellmath__62__W0[12], inst_cellmath__62__W0[11], inst_cellmath__62__W0[10], inst_cellmath__62__W0[9], inst_cellmath__62__W0[8], inst_cellmath__62__W0[7], inst_cellmath__62__W0[6], inst_cellmath__62__W0[5], inst_cellmath__62__W0[4], inst_cellmath__62__W0[3], inst_cellmath__62__W0[2], inst_cellmath__62__W0[1], inst_cellmath__62__W0[0]}));
cynw_cm_float_rcp_inst_cellmath__68_0_bdw1471647203_bdw cynw_cm_float_rcp_I31 (.inst_cellmath__68_0_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__68_0_in0(inst_cellmath__67), .inst_cellmath__68_0_in1({inst_cellmath__64[39], inst_cellmath__64[38], inst_cellmath__64[37], inst_cellmath__64[36], inst_cellmath__64[35], inst_cellmath__64[34], inst_cellmath__64[33], inst_cellmath__64[32], inst_cellmath__64[31], inst_cellmath__64[30], inst_cellmath__64[29], inst_cellmath__64[28], inst_cellmath__64[27], inst_cellmath__64[26], inst_cellmath__64[25], inst_cellmath__64[24], inst_cellmath__64[23], inst_cellmath__64[22], inst_cellmath__64[21], inst_cellmath__64[20], inst_cellmath__64[19], inst_cellmath__64[18], inst_cellmath__64[17]}), .inst_cellmath__68_0_in2(inst_cellmath__29));
assign inst_cellmath__19[1] = 1'B1;
assign inst_cellmath__19[2] = 1'B1;
assign inst_cellmath__19[3] = 1'B1;
assign inst_cellmath__19[4] = 1'B1;
assign inst_cellmath__19[5] = 1'B1;
assign inst_cellmath__19[6] = 1'B1;
assign inst_cellmath__19[7] = 1'B1;
assign inst_cellmath__19[8] = 1'B1;
assign inst_cellmath__48[0] = a_man[0];
assign inst_cellmath__48[1] = a_man[1];
assign inst_cellmath__48[2] = a_man[2];
assign inst_cellmath__48[3] = a_man[3];
assign inst_cellmath__48[4] = a_man[4];
assign inst_cellmath__48[5] = a_man[5];
assign inst_cellmath__48[6] = a_man[6];
assign inst_cellmath__48[7] = a_man[7];
assign inst_cellmath__48[8] = a_man[8];
assign inst_cellmath__48[9] = a_man[9];
assign inst_cellmath__48[10] = a_man[10];
assign inst_cellmath__48[11] = a_man[11];
assign inst_cellmath__48[12] = a_man[12];
assign inst_cellmath__48[13] = a_man[13];
assign inst_cellmath__48[14] = a_man[14];
assign inst_cellmath__51[18] = 1'B1;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_cellmath__9_0_bdw1471647203_bdw (
	inst_cellmath__9_0_out0,
	inst_cellmath__9_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__9_0_out0;
input [7:0] inst_cellmath__9_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2X1 inst_cellmath__9_0_I0 (.Y(N11), .A(inst_cellmath__9_0_in0[7]), .B(inst_cellmath__9_0_in0[0]));
NAND2XL inst_cellmath__9_0_I1 (.Y(N12), .A(inst_cellmath__9_0_in0[6]), .B(inst_cellmath__9_0_in0[5]));
NAND2X1 inst_cellmath__9_0_I2 (.Y(N13), .A(inst_cellmath__9_0_in0[4]), .B(inst_cellmath__9_0_in0[3]));
NAND2XL inst_cellmath__9_0_I3 (.Y(N14), .A(inst_cellmath__9_0_in0[2]), .B(inst_cellmath__9_0_in0[1]));
NOR2XL inst_cellmath__9_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__9_0_I5 (.Y(N16), .A(N13), .B(N14));
CLKAND2X2 inst_cellmath__9_0_I6 (.Y(inst_cellmath__9_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_rcp_inst_cellmath__15__5__bdw1471647203_bdw (
	inst_cellmath__15__5__out0,
	inst_cellmath__15__5__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__15__5__out0;
input [22:0] inst_cellmath__15__5__in0;
wire N26,N27,N28,N29,N30,N31,N32 
	,N33,N34,N35,N36,N37,N38,N39,N40 
	,N41,N42,N43,N44,N45,N47,N48;
NOR2XL inst_cellmath__15__5__I0 (.Y(N26), .A(inst_cellmath__15__5__in0[0]), .B(inst_cellmath__15__5__in0[1]));
NOR2XL inst_cellmath__15__5__I1 (.Y(N27), .A(inst_cellmath__15__5__in0[22]), .B(inst_cellmath__15__5__in0[21]));
NOR2XL inst_cellmath__15__5__I2 (.Y(N28), .A(inst_cellmath__15__5__in0[20]), .B(inst_cellmath__15__5__in0[19]));
NOR2XL inst_cellmath__15__5__I3 (.Y(N29), .A(inst_cellmath__15__5__in0[18]), .B(inst_cellmath__15__5__in0[17]));
NOR2XL inst_cellmath__15__5__I4 (.Y(N30), .A(inst_cellmath__15__5__in0[16]), .B(inst_cellmath__15__5__in0[15]));
NOR2XL inst_cellmath__15__5__I5 (.Y(N31), .A(inst_cellmath__15__5__in0[14]), .B(inst_cellmath__15__5__in0[13]));
NOR2XL inst_cellmath__15__5__I6 (.Y(N32), .A(inst_cellmath__15__5__in0[12]), .B(inst_cellmath__15__5__in0[11]));
NOR2XL inst_cellmath__15__5__I7 (.Y(N33), .A(inst_cellmath__15__5__in0[10]), .B(inst_cellmath__15__5__in0[9]));
NOR2XL inst_cellmath__15__5__I8 (.Y(N34), .A(inst_cellmath__15__5__in0[8]), .B(inst_cellmath__15__5__in0[7]));
NOR2XL inst_cellmath__15__5__I9 (.Y(N35), .A(inst_cellmath__15__5__in0[6]), .B(inst_cellmath__15__5__in0[5]));
NOR2XL inst_cellmath__15__5__I10 (.Y(N36), .A(inst_cellmath__15__5__in0[4]), .B(inst_cellmath__15__5__in0[3]));
INVXL inst_cellmath__15__5__I11 (.Y(N37), .A(inst_cellmath__15__5__in0[2]));
NAND2XL inst_cellmath__15__5__I12 (.Y(N38), .A(N37), .B(N26));
NAND2XL inst_cellmath__15__5__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__15__5__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__15__5__I15 (.Y(N41), .A(N31), .B(N32));
NAND2XL inst_cellmath__15__5__I16 (.Y(N42), .A(N33), .B(N34));
NAND2XL inst_cellmath__15__5__I17 (.Y(N43), .A(N35), .B(N36));
NOR2XL inst_cellmath__15__5__I18 (.Y(N44), .A(N38), .B(N39));
NOR2XL inst_cellmath__15__5__I19 (.Y(N45), .A(N40), .B(N41));
NAND2XL inst_cellmath__15__5__I21 (.Y(N47), .A(N44), .B(N45));
OR2XL inst_cellmath__15__5__I169 (.Y(N48), .A(N42), .B(N43));
NOR2XL inst_cellmath__15__5__I23 (.Y(inst_cellmath__15__5__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_rcp_inst_cellmath__29_0_bdw1471647203_bdw (
	inst_cellmath__29_0_out0,
	inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__29_0_out0;
input  inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1;
wire N5;
INVXL inst_cellmath__29_0_I0 (.Y(N5), .A(inst_cellmath__29_0_in0));
NOR2X1 inst_cellmath__29_0_I1 (.Y(inst_cellmath__29_0_out0), .A(N5), .B(inst_cellmath__29_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__37_0_bdw1471647203_bdw (
	inst_cellmath__37_0_out0,
	inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__37_0_out0;
input  inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1;
wire N5;
INVXL inst_cellmath__37_0_I0 (.Y(N5), .A(inst_cellmath__37_0_in1));
NOR2X1 inst_cellmath__37_0_I1 (.Y(inst_cellmath__37_0_out0), .A(N5), .B(inst_cellmath__37_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__28_0_bdw1471647203_bdw (
	inst_cellmath__28_0_out0,
	inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__28_0_out0;
input  inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1;
CLKAND2X2 inst_cellmath__28_0_I0 (.Y(inst_cellmath__28_0_out0), .A(inst_cellmath__28_0_in0), .B(inst_cellmath__28_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__22_0_bdw1471647203_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output [8:0] inst_cellmath__22_0_out0;
input [7:0] inst_cellmath__22_0_in0;
input  inst_cellmath__22_0_in1;
wire N63,N67,N73,N80,N84,N90,N102 
	,N149,N154,N159,N221,N239,N253,N261,N270 
	,N275,N276,N379;
CLKAND2X3 inst_cellmath__22_0_I19 (.Y(N63), .A(inst_cellmath__22_0_in0[0]), .B(inst_cellmath__22_0_in1));
INVXL inst_cellmath__22_0_I134 (.Y(N253), .A(N63));
NOR2X4 inst_cellmath__22_0_I23 (.Y(N67), .A(inst_cellmath__22_0_in0[1]), .B(N63));
NOR2XL inst_cellmath__22_0_I27 (.Y(N73), .A(inst_cellmath__22_0_in0[3]), .B(inst_cellmath__22_0_in0[2]));
INVXL inst_cellmath__22_0_I142 (.Y(N261), .A(N253));
NAND2BXL inst_cellmath__22_0_I266 (.Y(N80), .AN(inst_cellmath__22_0_in0[2]), .B(N67));
NAND2X4 inst_cellmath__22_0_I35 (.Y(N84), .A(N73), .B(N67));
NOR2XL inst_cellmath__22_0_I39 (.Y(N90), .A(inst_cellmath__22_0_in0[5]), .B(inst_cellmath__22_0_in0[4]));
INVXL inst_cellmath__22_0_I151 (.Y(N270), .A(inst_cellmath__22_0_in0[6]));
NAND2XL inst_cellmath__22_0_I49 (.Y(N102), .A(N270), .B(N90));
NOR3BXL inst_cellmath__22_0_I119 (.Y(N159), .AN(N90), .B(inst_cellmath__22_0_in0[7]), .C(inst_cellmath__22_0_in0[6]));
INVXL inst_cellmath__22_0_I156 (.Y(N275), .A(inst_cellmath__22_0_in0[5]));
INVXL inst_cellmath__22_0_I157 (.Y(N276), .A(inst_cellmath__22_0_in0[7]));
XOR2XL inst_cellmath__22_0_I77 (.Y(inst_cellmath__22_0_out0[0]), .A(inst_cellmath__22_0_in0[0]), .B(inst_cellmath__22_0_in1));
INVXL xnor2_A_I106 (.Y(N221), .A(N261));
MXI2X1 xnor2_A_I107 (.Y(inst_cellmath__22_0_out0[1]), .A(N261), .B(N221), .S0(inst_cellmath__22_0_in0[1]));
XOR2XL inst_cellmath__22_0_I275 (.Y(inst_cellmath__22_0_out0[2]), .A(N67), .B(inst_cellmath__22_0_in0[2]));
XNOR2X1 inst_cellmath__22_0_I269 (.Y(inst_cellmath__22_0_out0[3]), .A(N80), .B(inst_cellmath__22_0_in0[3]));
INVXL xnor2_A_I112 (.Y(N239), .A(N84));
MXI2XL xnor2_A_I113 (.Y(inst_cellmath__22_0_out0[4]), .A(N84), .B(N239), .S0(inst_cellmath__22_0_in0[4]));
NOR2XL node_cs_const1_cs_A_I283 (.Y(N379), .A(inst_cellmath__22_0_in0[4]), .B(N84));
XNOR2X1 node_cs_const1_cs_A_I284 (.Y(inst_cellmath__22_0_out0[5]), .A(N275), .B(N379));
XOR2XL inst_cellmath__22_0_I173 (.Y(N149), .A(N90), .B(N270));
MXI2XL inst_cellmath__22_0_I85 (.Y(inst_cellmath__22_0_out0[6]), .A(N149), .B(N270), .S0(N84));
XNOR2X1 inst_cellmath__22_0_I86 (.Y(N154), .A(N102), .B(N276));
MXI2XL inst_cellmath__22_0_I87 (.Y(inst_cellmath__22_0_out0[7]), .A(N154), .B(N276), .S0(N84));
NOR2BXL inst_cellmath__22_0_I273 (.Y(inst_cellmath__22_0_out0[8]), .AN(N159), .B(N84));
endmodule

module cynw_cm_float_rcp_inst_cellmath__17__6__bdw1471647203_bdw (
	inst_cellmath__17__6__out0,
	inst_cellmath__17__6__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__17__6__out0;
input [7:0] inst_cellmath__17__6__in0;
wire N17,N18,N19,N20;
NOR3X1 inst_cellmath__17__6__I13 (.Y(N18), .A(inst_cellmath__17__6__in0[0]), .B(inst_cellmath__17__6__in0[1]), .C(inst_cellmath__17__6__in0[4]));
NOR3XL inst_cellmath__17__6__I26 (.Y(N20), .A(inst_cellmath__17__6__in0[2]), .B(inst_cellmath__17__6__in0[3]), .C(inst_cellmath__17__6__in0[5]));
NOR2X2 inst_cellmath__17__6__I6 (.Y(N17), .A(inst_cellmath__17__6__in0[6]), .B(inst_cellmath__17__6__in0[7]));
CLKAND2X3 inst_cellmath__17__6__I8 (.Y(N19), .A(N18), .B(N17));
NAND2X1 inst_cellmath__17__6__I10 (.Y(inst_cellmath__17__6__out0[0]), .A(N20), .B(N19));
endmodule

module cynw_cm_float_rcp_inst_cellmath__17_0_bdw1471647203_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0,
	inst_cellmath__17_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [8:8] inst_cellmath__17_0_in0;
input [0:0] inst_cellmath__17_0_in1;
NAND2BX2 inst_cellmath__17_0_I4 (.Y(inst_cellmath__17_0_out0), .AN(inst_cellmath__17_0_in0[8]), .B(inst_cellmath__17_0_in1[0]));
endmodule

module cynw_cm_float_rcp_inst_cellmath__30_0_bdw1471647203_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__30_0_out0;
input  inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
wire N5;
INVXL inst_cellmath__30_0_I0 (.Y(N5), .A(inst_cellmath__30_0_in0));
CLKAND2X6 inst_cellmath__30_0_I1 (.Y(inst_cellmath__30_0_out0), .A(N5), .B(inst_cellmath__30_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__33__7__bdw1471647203_bdw (
	inst_cellmath__33__7__out0,
	inst_cellmath__33__7__in0,
	inst_cellmath__33__7__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__33__7__out0;
input  inst_cellmath__33__7__in0,
	inst_cellmath__33__7__in1;
OR2XL inst_cellmath__33__7__I0 (.Y(inst_cellmath__33__7__out0[0]), .A(inst_cellmath__33__7__in1), .B(inst_cellmath__33__7__in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__33_0_bdw1471647203_bdw (
	inst_cellmath__33_0_out0,
	inst_cellmath__33_0_in0,
	inst_cellmath__33_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__33_0_out0;
input [0:0] inst_cellmath__33_0_in0;
input  inst_cellmath__33_0_in1;
wire N5;
INVXL inst_cellmath__33_0_I0 (.Y(N5), .A(inst_cellmath__33_0_in1));
CLKAND2X6 inst_cellmath__33_0_I1 (.Y(inst_cellmath__33_0_out0), .A(N5), .B(inst_cellmath__33_0_in0[0]));
endmodule

module cynw_cm_float_rcp_inst_cellmath__34_0_bdw1471647203_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0,
	inst_cellmath__34_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__34_0_out0;
input  inst_cellmath__34_0_in0;
input [7:0] inst_cellmath__34_0_in1;
wire N12,N13,N14,N15,N19;
NOR2XL inst_cellmath__34_0_I0 (.Y(N12), .A(inst_cellmath__34_0_in1[0]), .B(inst_cellmath__34_0_in1[1]));
NOR2XL inst_cellmath__34_0_I1 (.Y(N13), .A(inst_cellmath__34_0_in1[7]), .B(inst_cellmath__34_0_in1[6]));
NOR2XL inst_cellmath__34_0_I2 (.Y(N14), .A(inst_cellmath__34_0_in1[5]), .B(inst_cellmath__34_0_in1[4]));
NOR2XL inst_cellmath__34_0_I3 (.Y(N15), .A(inst_cellmath__34_0_in1[3]), .B(inst_cellmath__34_0_in1[2]));
NAND4XL inst_cellmath__34_0_I11 (.Y(N19), .A(N12), .B(N14), .C(N13), .D(N15));
NOR2X1 inst_cellmath__34_0_I8 (.Y(inst_cellmath__34_0_out0), .A(N19), .B(inst_cellmath__34_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__42__9__bdw1471647203_bdw (
	inst_cellmath__42__9__out0,
	inst_cellmath__42__9__in0,
	inst_cellmath__42__9__in1,
	inst_cellmath__42__9__in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__42__9__out0;
input  inst_cellmath__42__9__in0,
	inst_cellmath__42__9__in1,
	inst_cellmath__42__9__in2;
wire N7;
OR2XL inst_cellmath__42__9__I0 (.Y(N7), .A(inst_cellmath__42__9__in2), .B(inst_cellmath__42__9__in0));
NOR2X2 inst_cellmath__42__9__I2 (.Y(inst_cellmath__42__9__out0), .A(N7), .B(inst_cellmath__42__9__in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__38_0_bdw1471647203_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1;
OR2XL inst_cellmath__38_0_I0 (.Y(inst_cellmath__38_0_out0), .A(inst_cellmath__38_0_in1), .B(inst_cellmath__38_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__43_0_bdw1471647203_bdw (
	inst_cellmath__43_0_out0,
	inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1,
	inst_cellmath__43_0_in2
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__43_0_out0;
input  inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1;
input [7:0] inst_cellmath__43_0_in2;
MX2XL inst_cellmath__43_0_I16 (.Y(inst_cellmath__43_0_out0[0]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[0]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I17 (.Y(inst_cellmath__43_0_out0[1]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[1]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I18 (.Y(inst_cellmath__43_0_out0[2]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[2]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I19 (.Y(inst_cellmath__43_0_out0[3]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[3]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I20 (.Y(inst_cellmath__43_0_out0[4]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[4]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I21 (.Y(inst_cellmath__43_0_out0[5]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[5]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I22 (.Y(inst_cellmath__43_0_out0[6]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[6]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I23 (.Y(inst_cellmath__43_0_out0[7]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[7]), .S0(inst_cellmath__43_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__67__11__bdw1471647203_bdw (
	inst_cellmath__67__11__out0,
	inst_cellmath__67__11__in0,
	inst_cellmath__67__11__in1,
	inst_cellmath__67__11__in2,
	inst_cellmath__67__11__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__67__11__out0;
input  inst_cellmath__67__11__in0,
	inst_cellmath__67__11__in1,
	inst_cellmath__67__11__in2,
	inst_cellmath__67__11__in3;
wire N10;
OR3XL inst_cellmath__67__11__I7 (.Y(N10), .A(inst_cellmath__67__11__in3), .B(inst_cellmath__67__11__in2), .C(inst_cellmath__67__11__in0));
OR2XL inst_cellmath__67__11__I4 (.Y(inst_cellmath__67__11__out0[0]), .A(N10), .B(inst_cellmath__67__11__in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__60_0_bdw1471647203_bdw (
	inst_cellmath__60_0_out0,
	inst_cellmath__60_0_in0,
	inst_cellmath__60_0_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__60_0_out0;
input  inst_cellmath__60_0_in0;
input [14:3] inst_cellmath__60_0_in1;
wire N80,N84,N86,N88,N90,N92,N94 
	,N96,N98,N100,N118,N120,N122,N124,N126 
	,N128,N130,N132,N134,N136,N150,N154,N156 
	,N158,N160,N162,N164,N166,N168,N170,N184 
	,N188,N190,N192,N194,N196,N198,N200,N202 
	,N216,N220,N222,N224,N226,N228,N230,N232 
	,N246,N250,N252,N254,N256,N258,N260,N274 
	,N278,N280,N282,N284,N286,N300,N304,N306 
	,N308,N310,N324,N328,N330,N332,N346,N350 
	,N352,N366,N370,N384,N404,N405,N406,N407 
	,N408,N409,N410,N411,N412,N413,N414,N415 
	,N416,N417,N418,N419,N420,N421,N422,N423 
	,N424,N425,N426,N427,N428,N429,N430,N431 
	,N432,N433,N434,N435,N436,N437,N438,N439 
	,N440,N441,N442,N443,N444,N445,N446,N447 
	,N448,N449,N450,N451,N452,N453,N454,N455 
	,N456,N457,N458,N459,N460,N461,N462,N463 
	,N464,N465,N466,N469,N470,N471,N472,N473 
	,N474,N475,N476,N477,N478,N479,N480,N481 
	,N482,N483,N484,N485,N486,N487,N488,N489 
	,N490,N491,N492,N493,N494,N495,N496,N497 
	,N498,N499,N500,N501,N502,N503,N504,N505 
	,N506,N507,N508,N509,N510,N511,N512,N513 
	,N514,N515,N516,N517,N518,N519,N520,N521 
	,N522,N523,N524,N525,N526,N527,N528,N529 
	,N530,N531,N532,N533,N534,N535,N536,N537 
	,N538,N539,N540,N543,N553,N561,N573,N585 
	,N601,N636,N639,N642,N645,N648,N651,N660 
	,N662,N663,N664,N665,N666,N667,N668,N669 
	,N670,N671,N672,N673,N674,N675,N676,N677 
	,N678,N679,N680,N681,N682,N683,N684,N685 
	,N686,N687,N688,N689,N694,N698,N699,N702 
	,N703,N706,N707,N710,N711,N714,N715,N718 
	,N719,N724,N742,N744,N745,N746,N747,N748 
	,N749,N750,N751,N756,N758,N760,N761,N762 
	,N763,N772,N774,N801,N804,N807,N810,N813 
	,N816,N819,N822,N825,N828,N831,N834,N837 
	,N840,N843,N852,N853,N855,N856,N858,N859 
	,N861,N862,N864,N865,N867,N868,N870,N871 
	,N873,N874,N1057,N1066,N1109,N1111,N1115,N1119 
	,N1124,N1126,N1127,N1128,N1131,N1133,N1137,N1138 
	,N1143,N1148,N1153,N1158,N1161,N1162,N1168,N1169 
	,N1179,N1180,N1206,N1207,N1220,N1221,N1222,N1223 
	,N1224,N1241,N1253,N1260;
INVXL inst_cellmath__60_0_I654 (.Y(N1111), .A(inst_cellmath__60_0_in1[4]));
INVX1 inst_cellmath__60_0_I652 (.Y(N1109), .A(inst_cellmath__60_0_in1[4]));
INVX2 inst_cellmath__60_0_I658 (.Y(N1115), .A(inst_cellmath__60_0_in1[5]));
INVX2 inst_cellmath__60_0_I662 (.Y(N1119), .A(inst_cellmath__60_0_in1[6]));
INVX3 inst_cellmath__60_0_I667 (.Y(N1124), .A(inst_cellmath__60_0_in1[7]));
INVX2 inst_cellmath__60_0_I669 (.Y(N1126), .A(inst_cellmath__60_0_in1[8]));
INVX2 inst_cellmath__60_0_I670 (.Y(N1127), .A(inst_cellmath__60_0_in1[9]));
INVX2 inst_cellmath__60_0_I671 (.Y(N1128), .A(inst_cellmath__60_0_in1[10]));
INVX1 inst_cellmath__60_0_I676 (.Y(N1133), .A(inst_cellmath__60_0_in1[11]));
INVXL inst_cellmath__60_0_I674 (.Y(N1131), .A(inst_cellmath__60_0_in1[11]));
INVXL inst_cellmath__60_0_I681 (.Y(N1138), .A(inst_cellmath__60_0_in1[12]));
INVX1 inst_cellmath__60_0_I680 (.Y(N1137), .A(inst_cellmath__60_0_in1[12]));
INVX2 inst_cellmath__60_0_I686 (.Y(N1143), .A(inst_cellmath__60_0_in1[13]));
INVX2 inst_cellmath__60_0_I691 (.Y(N1148), .A(inst_cellmath__60_0_in1[14]));
INVX1 inst_cellmath__60_0_I696 (.Y(N1153), .A(inst_cellmath__60_0_in0));
INVX2 inst_cellmath__60_0_I701 (.Y(N1158), .A(inst_cellmath__60_0_in1[3]));
INVXL inst_cellmath__60_0_I17 (.Y(inst_cellmath__60_0_out0[0]), .A(N1158));
OR2XL inst_cellmath__60_0_I19 (.Y(N80), .A(N1158), .B(N1111));
NOR2XL inst_cellmath__60_0_I20 (.Y(N528), .A(N1158), .B(N1115));
NOR2BX1 inst_cellmath__60_0_I801 (.Y(N84), .AN(inst_cellmath__60_0_in1[6]), .B(N1158));
NOR2BX1 inst_cellmath__60_0_I802 (.Y(N86), .AN(inst_cellmath__60_0_in1[7]), .B(N1158));
NOR2XL inst_cellmath__60_0_I23 (.Y(N88), .A(N1158), .B(N1126));
NOR2XL inst_cellmath__60_0_I24 (.Y(N90), .A(N1158), .B(N1127));
NOR2XL inst_cellmath__60_0_I25 (.Y(N92), .A(N1158), .B(N1128));
NOR2XL inst_cellmath__60_0_I26 (.Y(N94), .A(N1158), .B(N1133));
NOR2XL inst_cellmath__60_0_I27 (.Y(N96), .A(N1158), .B(N1138));
NOR2XL inst_cellmath__60_0_I28 (.Y(N98), .A(N1158), .B(N1143));
NOR2XL inst_cellmath__60_0_I29 (.Y(N100), .A(N1158), .B(N1148));
OR2XL inst_cellmath__60_0_I30 (.Y(N404), .A(N1158), .B(N1153));
NOR2XL inst_cellmath__60_0_I37 (.Y(N118), .A(N1111), .B(N1115));
NOR2XL inst_cellmath__60_0_I38 (.Y(N120), .A(N1111), .B(N1119));
NOR2XL inst_cellmath__60_0_I39 (.Y(N122), .A(N1111), .B(N1124));
NOR2XL inst_cellmath__60_0_I40 (.Y(N124), .A(N1111), .B(N1126));
NOR2XL inst_cellmath__60_0_I41 (.Y(N126), .A(N1111), .B(N1127));
NOR2XL inst_cellmath__60_0_I42 (.Y(N128), .A(N1111), .B(N1128));
NOR2XL inst_cellmath__60_0_I43 (.Y(N130), .A(N1109), .B(N1133));
NOR2XL inst_cellmath__60_0_I44 (.Y(N132), .A(N1109), .B(N1138));
NOR2X1 inst_cellmath__60_0_I45 (.Y(N134), .A(N1109), .B(N1143));
NOR2XL inst_cellmath__60_0_I46 (.Y(N136), .A(N1109), .B(N1148));
OR2XL inst_cellmath__60_0_I47 (.Y(N405), .A(N1109), .B(N1153));
INVXL inst_cellmath__60_0_I52 (.Y(N150), .A(N1115));
NOR2XL inst_cellmath__60_0_I54 (.Y(N154), .A(N1115), .B(N1119));
NOR2XL inst_cellmath__60_0_I55 (.Y(N156), .A(N1115), .B(N1124));
NOR2XL inst_cellmath__60_0_I56 (.Y(N158), .A(N1115), .B(N1126));
NOR2XL inst_cellmath__60_0_I57 (.Y(N160), .A(N1115), .B(N1127));
NOR2XL inst_cellmath__60_0_I58 (.Y(N162), .A(N1115), .B(N1128));
NOR2XL inst_cellmath__60_0_I59 (.Y(N164), .A(N1115), .B(N1133));
NOR2XL inst_cellmath__60_0_I60 (.Y(N166), .A(N1115), .B(N1138));
NOR2XL inst_cellmath__60_0_I61 (.Y(N168), .A(N1115), .B(N1143));
NOR2XL inst_cellmath__60_0_I62 (.Y(N170), .A(N1115), .B(N1148));
OR2XL inst_cellmath__60_0_I63 (.Y(N406), .A(N1115), .B(N1153));
INVXL inst_cellmath__60_0_I68 (.Y(N184), .A(N1119));
NOR2XL inst_cellmath__60_0_I70 (.Y(N188), .A(N1119), .B(N1124));
NOR2XL inst_cellmath__60_0_I71 (.Y(N190), .A(N1119), .B(N1126));
NOR2XL inst_cellmath__60_0_I72 (.Y(N192), .A(N1119), .B(N1127));
NOR2XL inst_cellmath__60_0_I73 (.Y(N194), .A(N1119), .B(N1128));
NOR2XL inst_cellmath__60_0_I74 (.Y(N196), .A(N1119), .B(N1133));
NOR2X1 inst_cellmath__60_0_I75 (.Y(N198), .A(N1119), .B(N1137));
NOR2XL inst_cellmath__60_0_I76 (.Y(N200), .A(N1119), .B(N1143));
NOR2XL inst_cellmath__60_0_I77 (.Y(N202), .A(N1119), .B(N1148));
OR2XL inst_cellmath__60_0_I78 (.Y(N407), .A(N1119), .B(N1153));
INVXL inst_cellmath__60_0_I83 (.Y(N216), .A(N1124));
NOR2XL inst_cellmath__60_0_I85 (.Y(N220), .A(N1124), .B(N1126));
NOR2XL inst_cellmath__60_0_I86 (.Y(N222), .A(N1124), .B(N1127));
NOR2X2 inst_cellmath__60_0_I87 (.Y(N224), .A(N1124), .B(N1128));
NOR2X1 inst_cellmath__60_0_I88 (.Y(N226), .A(N1124), .B(N1133));
NOR2X1 inst_cellmath__60_0_I89 (.Y(N228), .A(N1124), .B(N1137));
NOR2XL inst_cellmath__60_0_I90 (.Y(N230), .A(N1124), .B(N1143));
NOR2XL inst_cellmath__60_0_I91 (.Y(N232), .A(N1124), .B(N1148));
OR2XL inst_cellmath__60_0_I92 (.Y(N408), .A(N1124), .B(N1153));
INVXL inst_cellmath__60_0_I97 (.Y(N246), .A(N1126));
NOR2X2 inst_cellmath__60_0_I99 (.Y(N250), .A(N1126), .B(N1127));
NOR2XL inst_cellmath__60_0_I100 (.Y(N252), .A(N1126), .B(N1128));
NOR2X1 inst_cellmath__60_0_I101 (.Y(N254), .A(N1126), .B(N1133));
NOR2XL inst_cellmath__60_0_I102 (.Y(N256), .A(N1126), .B(N1137));
NOR2X1 inst_cellmath__60_0_I103 (.Y(N258), .A(N1126), .B(N1143));
NOR2XL inst_cellmath__60_0_I104 (.Y(N260), .A(N1126), .B(N1148));
OR2XL inst_cellmath__60_0_I105 (.Y(N409), .A(N1126), .B(N1153));
INVXL inst_cellmath__60_0_I110 (.Y(N274), .A(N1127));
NOR2X1 inst_cellmath__60_0_I112 (.Y(N278), .A(N1127), .B(N1128));
NOR2XL inst_cellmath__60_0_I113 (.Y(N280), .A(N1127), .B(N1133));
NOR2XL inst_cellmath__60_0_I114 (.Y(N282), .A(N1127), .B(N1137));
NOR2XL inst_cellmath__60_0_I115 (.Y(N284), .A(N1127), .B(N1143));
NOR2XL inst_cellmath__60_0_I116 (.Y(N286), .A(N1127), .B(N1148));
OR2XL inst_cellmath__60_0_I117 (.Y(N410), .A(N1127), .B(N1153));
INVXL inst_cellmath__60_0_I122 (.Y(N300), .A(N1128));
NOR2X1 inst_cellmath__60_0_I124 (.Y(N304), .A(N1128), .B(N1133));
NOR2XL inst_cellmath__60_0_I125 (.Y(N306), .A(N1128), .B(N1137));
NOR2XL inst_cellmath__60_0_I126 (.Y(N308), .A(N1128), .B(N1143));
NOR2XL inst_cellmath__60_0_I127 (.Y(N310), .A(N1128), .B(N1148));
OR2XL inst_cellmath__60_0_I128 (.Y(N411), .A(N1128), .B(N1153));
INVXL inst_cellmath__60_0_I133 (.Y(N324), .A(N1131));
NOR2XL inst_cellmath__60_0_I135 (.Y(N328), .A(N1131), .B(N1138));
NOR2XL inst_cellmath__60_0_I136 (.Y(N330), .A(N1131), .B(N1143));
NOR2XL inst_cellmath__60_0_I137 (.Y(N332), .A(N1131), .B(N1148));
OR2XL inst_cellmath__60_0_I138 (.Y(N412), .A(N1131), .B(N1153));
INVXL inst_cellmath__60_0_I143 (.Y(N346), .A(N1138));
NOR2XL inst_cellmath__60_0_I145 (.Y(N350), .A(N1138), .B(N1143));
NOR2XL inst_cellmath__60_0_I146 (.Y(N352), .A(N1138), .B(N1148));
OR2XL inst_cellmath__60_0_I147 (.Y(N413), .A(N1138), .B(N1153));
INVXL inst_cellmath__60_0_I152 (.Y(N366), .A(N1143));
NOR2XL inst_cellmath__60_0_I154 (.Y(N370), .A(N1143), .B(N1148));
OR2XL inst_cellmath__60_0_I155 (.Y(N414), .A(N1143), .B(N1153));
INVXL inst_cellmath__60_0_I160 (.Y(N384), .A(N1148));
ADDHX1 inst_cellmath__60_0_I179 (.CO(N416), .S(N415), .A(N150), .B(N84));
ADDHX1 inst_cellmath__60_0_I180 (.CO(N418), .S(N417), .A(N120), .B(N86));
ADDHX1 inst_cellmath__60_0_I181 (.CO(N420), .S(N419), .A(N184), .B(N88));
ADDFX1 inst_cellmath__60_0_I182 (.CO(N422), .S(N421), .A(N154), .B(N122), .CI(N418));
ADDHX1 inst_cellmath__60_0_I183 (.CO(N424), .S(N423), .A(N156), .B(N90));
ADDFX1 inst_cellmath__60_0_I184 (.CO(N426), .S(N425), .A(N420), .B(N124), .CI(N423));
ADDHX1 inst_cellmath__60_0_I185 (.CO(N428), .S(N427), .A(N216), .B(N92));
ADDFX1 inst_cellmath__60_0_I186 (.CO(N430), .S(N429), .A(N158), .B(N188), .CI(N126));
ADDFX1 inst_cellmath__60_0_I187 (.CO(N432), .S(N431), .A(N427), .B(N424), .CI(N429));
ADDHX1 inst_cellmath__60_0_I188 (.CO(N434), .S(N433), .A(N190), .B(N94));
ADDFX1 inst_cellmath__60_0_I189 (.CO(N436), .S(N435), .A(N128), .B(N160), .CI(N428));
ADDFX1 inst_cellmath__60_0_I190 (.CO(N438), .S(N437), .A(N430), .B(N433), .CI(N435));
ADDHX1 inst_cellmath__60_0_I191 (.CO(N440), .S(N439), .A(N246), .B(N96));
ADDFX1 inst_cellmath__60_0_I192 (.CO(N442), .S(N441), .A(N192), .B(N220), .CI(N130));
ADDFX1 inst_cellmath__60_0_I193 (.CO(N444), .S(N443), .A(N434), .B(N162), .CI(N439));
ADDFX1 inst_cellmath__60_0_I194 (.CO(N446), .S(N445), .A(N436), .B(N441), .CI(N443));
ADDHX1 inst_cellmath__60_0_I195 (.CO(N448), .S(N447), .A(N222), .B(N98));
ADDFX1 inst_cellmath__60_0_I196 (.CO(N450), .S(N449), .A(N164), .B(N194), .CI(N132));
ADDFX1 inst_cellmath__60_0_I197 (.CO(N452), .S(N451), .A(N447), .B(N440), .CI(N442));
ADDFX1 inst_cellmath__60_0_I198 (.CO(N454), .S(N453), .A(N444), .B(N449), .CI(N451));
ADDHX1 inst_cellmath__60_0_I199 (.CO(N456), .S(N455), .A(N274), .B(N100));
ADDFX1 inst_cellmath__60_0_I200 (.CO(N458), .S(N457), .A(N224), .B(N250), .CI(N134));
ADDFX1 inst_cellmath__60_0_I201 (.CO(N460), .S(N459), .A(N166), .B(N196), .CI(N448));
ADDFX1 inst_cellmath__60_0_I202 (.CO(N462), .S(N461), .A(N450), .B(N455), .CI(N457));
ADDFX1 inst_cellmath__60_0_I203 (.CO(N464), .S(N463), .A(N452), .B(N459), .CI(N461));
XNOR2X1 hap1_A_I598 (.Y(N465), .A(N252), .B(N168));
OR2XL hap1_A_I599 (.Y(N466), .A(N252), .B(N168));
ADDFX1 inst_cellmath__60_0_I205 (.CO(N470), .S(N469), .A(N198), .B(N226), .CI(N136));
ADDFHXL inst_cellmath__60_0_I206 (.CO(N472), .S(N471), .A(N456), .B(N404), .CI(N458));
ADDFX1 inst_cellmath__60_0_I207 (.CO(N474), .S(N473), .A(N469), .B(N465), .CI(N460));
ADDFX1 inst_cellmath__60_0_I208 (.CO(N476), .S(N475), .A(N462), .B(N471), .CI(N473));
ADDFX1 inst_cellmath__60_0_I209 (.CO(N478), .S(N477), .A(N278), .B(N300), .CI(N200));
ADDFX1 inst_cellmath__60_0_I210 (.CO(N480), .S(N479), .A(N228), .B(N254), .CI(N170));
ADDFX1 inst_cellmath__60_0_I211 (.CO(N482), .S(N481), .A(N466), .B(N405), .CI(N470));
ADDFHXL inst_cellmath__60_0_I212 (.CO(N484), .S(N483), .A(N479), .B(N477), .CI(N472));
ADDFHX1 inst_cellmath__60_0_I213 (.CO(N486), .S(N485), .A(N474), .B(N481), .CI(N483));
ADDFX1 inst_cellmath__60_0_I214 (.CO(N488), .S(N487), .A(N256), .B(N280), .CI(N202));
ADDFX1 inst_cellmath__60_0_I215 (.CO(N490), .S(N489), .A(N406), .B(N230), .CI(N478));
ADDFXL inst_cellmath__60_0_I216 (.CO(N492), .S(N491), .A(N487), .B(N480), .CI(N482));
ADDFX1 inst_cellmath__60_0_I217 (.CO(N494), .S(N493), .A(N484), .B(N489), .CI(N491));
ADDFX1 inst_cellmath__60_0_I218 (.CO(N496), .S(N495), .A(N304), .B(N324), .CI(N232));
ADDFX1 inst_cellmath__60_0_I219 (.CO(N498), .S(N497), .A(N258), .B(N282), .CI(N407));
ADDFXL inst_cellmath__60_0_I220 (.CO(N500), .S(N499), .A(N495), .B(N488), .CI(N497));
ADDFHX1 inst_cellmath__60_0_I221 (.CO(N502), .S(N501), .A(N492), .B(N490), .CI(N499));
ADDFX1 inst_cellmath__60_0_I222 (.CO(N504), .S(N503), .A(N284), .B(N306), .CI(N260));
ADDFX1 inst_cellmath__60_0_I223 (.CO(N506), .S(N505), .A(N496), .B(N408), .CI(N498));
ADDFX1 inst_cellmath__60_0_I224 (.CO(N508), .S(N507), .A(N500), .B(N503), .CI(N505));
ADDFX1 inst_cellmath__60_0_I225 (.CO(N510), .S(N509), .A(N328), .B(N346), .CI(N286));
ADDFX1 inst_cellmath__60_0_I226 (.CO(N512), .S(N511), .A(N409), .B(N308), .CI(N504));
ADDFX1 inst_cellmath__60_0_I227 (.CO(N514), .S(N513), .A(N506), .B(N509), .CI(N511));
ADDFX1 inst_cellmath__60_0_I228 (.CO(N516), .S(N515), .A(N310), .B(N330), .CI(N410));
ADDFX1 inst_cellmath__60_0_I229 (.CO(N518), .S(N517), .A(N515), .B(N510), .CI(N512));
ADDFX1 inst_cellmath__60_0_I230 (.CO(N520), .S(N519), .A(N350), .B(N366), .CI(N332));
ADDFX1 inst_cellmath__60_0_I231 (.CO(N522), .S(N521), .A(N516), .B(N411), .CI(N519));
ADDFX1 inst_cellmath__60_0_I232 (.CO(N524), .S(N523), .A(N412), .B(N352), .CI(N520));
ADDFX1 inst_cellmath__60_0_I233 (.CO(N526), .S(N525), .A(N370), .B(N384), .CI(N413));
NOR2XL inst_cellmath__60_0_I234 (.Y(N527), .A(N1109), .B(N80));
NOR2XL inst_cellmath__60_0_I236 (.Y(N529), .A(N118), .B(N415));
NAND2XL inst_cellmath__60_0_I237 (.Y(N530), .A(N118), .B(N415));
NOR2XL inst_cellmath__60_0_I238 (.Y(N531), .A(N416), .B(N417));
NAND2XL inst_cellmath__60_0_I239 (.Y(N532), .A(N416), .B(N417));
NOR2XL inst_cellmath__60_0_I240 (.Y(N533), .A(N419), .B(N421));
NAND2XL inst_cellmath__60_0_I241 (.Y(N534), .A(N419), .B(N421));
NOR2XL inst_cellmath__60_0_I242 (.Y(N535), .A(N422), .B(N425));
NAND2XL inst_cellmath__60_0_I243 (.Y(N536), .A(N422), .B(N425));
NOR2XL inst_cellmath__60_0_I244 (.Y(N537), .A(N426), .B(N431));
NAND2XL inst_cellmath__60_0_I245 (.Y(N538), .A(N426), .B(N431));
NOR2XL inst_cellmath__60_0_I246 (.Y(N539), .A(N432), .B(N437));
NAND2XL inst_cellmath__60_0_I247 (.Y(N540), .A(N432), .B(N437));
AND2XL inst_cellmath__60_0_I250 (.Y(N543), .A(N528), .B(N527));
INVXL inst_cellmath__60_0_I704 (.Y(N1161), .A(N529));
INVXL inst_cellmath__60_0_I705 (.Y(N1162), .A(N530));
OAI21XL inst_cellmath__60_0_I258 (.Y(N553), .A0(N1162), .A1(N543), .B0(N1161));
AOI21XL inst_cellmath__60_0_I266 (.Y(N561), .A0(N532), .A1(N553), .B0(N531));
INVXL inst_cellmath__60_0_I711 (.Y(N1168), .A(N533));
INVXL inst_cellmath__60_0_I712 (.Y(N1169), .A(N534));
OAI21X2 inst_cellmath__60_0_I278 (.Y(N573), .A0(N1169), .A1(N561), .B0(N1168));
AOI21X2 inst_cellmath__60_0_I290 (.Y(N585), .A0(N536), .A1(N573), .B0(N535));
INVXL inst_cellmath__60_0_I722 (.Y(N1179), .A(N537));
INVXL inst_cellmath__60_0_I723 (.Y(N1180), .A(N538));
OAI21X1 inst_cellmath__60_0_I306 (.Y(N601), .A0(N1180), .A1(N585), .B0(N1179));
NAND2BXL inst_cellmath__60_0_I339 (.Y(N636), .AN(N529), .B(N530));
NAND2BXL inst_cellmath__60_0_I342 (.Y(N639), .AN(N531), .B(N532));
NAND2BXL inst_cellmath__60_0_I345 (.Y(N642), .AN(N533), .B(N534));
NAND2BXL inst_cellmath__60_0_I348 (.Y(N645), .AN(N535), .B(N536));
NAND2BXL inst_cellmath__60_0_I351 (.Y(N648), .AN(N537), .B(N538));
NAND2BXL inst_cellmath__60_0_I354 (.Y(N651), .AN(N539), .B(N540));
XOR2XL inst_cellmath__60_0_I355 (.Y(inst_cellmath__60_0_out0[2]), .A(N1111), .B(N80));
XOR2XL inst_cellmath__60_0_I803 (.Y(inst_cellmath__60_0_out0[3]), .A(N527), .B(N528));
XNOR2X1 inst_cellmath__60_0_I357 (.Y(inst_cellmath__60_0_out0[4]), .A(N543), .B(N636));
XOR2XL inst_cellmath__60_0_I804 (.Y(inst_cellmath__60_0_out0[5]), .A(N553), .B(N639));
XNOR2X1 inst_cellmath__60_0_I359 (.Y(inst_cellmath__60_0_out0[6]), .A(N561), .B(N642));
XOR2XL inst_cellmath__60_0_I805 (.Y(inst_cellmath__60_0_out0[7]), .A(N573), .B(N645));
XNOR2X1 inst_cellmath__60_0_I361 (.Y(inst_cellmath__60_0_out0[8]), .A(N585), .B(N648));
XOR2XL inst_cellmath__60_0_I806 (.Y(inst_cellmath__60_0_out0[9]), .A(N601), .B(N651));
AO21XL inst_cellmath__60_0_I857 (.Y(N660), .A0(N540), .A1(N601), .B0(N539));
NOR2XL inst_cellmath__60_0_I364 (.Y(N662), .A(N438), .B(N445));
NAND2XL inst_cellmath__60_0_I365 (.Y(N663), .A(N438), .B(N445));
NOR2X1 inst_cellmath__60_0_I366 (.Y(N664), .A(N446), .B(N453));
NAND2XL inst_cellmath__60_0_I367 (.Y(N665), .A(N446), .B(N453));
NOR2X1 inst_cellmath__60_0_I368 (.Y(N666), .A(N454), .B(N463));
NAND2X2 inst_cellmath__60_0_I369 (.Y(N667), .A(N454), .B(N463));
NOR2X2 inst_cellmath__60_0_I370 (.Y(N668), .A(N464), .B(N475));
NAND2X2 inst_cellmath__60_0_I371 (.Y(N669), .A(N464), .B(N475));
NOR2X1 inst_cellmath__60_0_I372 (.Y(N670), .A(N476), .B(N485));
NAND2X6 inst_cellmath__60_0_I373 (.Y(N671), .A(N476), .B(N485));
NOR2X2 inst_cellmath__60_0_I374 (.Y(N672), .A(N486), .B(N493));
NAND2X2 inst_cellmath__60_0_I375 (.Y(N673), .A(N486), .B(N493));
NOR2X1 inst_cellmath__60_0_I376 (.Y(N674), .A(N494), .B(N501));
NAND2X4 inst_cellmath__60_0_I377 (.Y(N675), .A(N494), .B(N501));
NOR2XL inst_cellmath__60_0_I378 (.Y(N676), .A(N502), .B(N507));
NAND2X1 inst_cellmath__60_0_I379 (.Y(N677), .A(N502), .B(N507));
NOR2XL inst_cellmath__60_0_I380 (.Y(N678), .A(N508), .B(N513));
NAND2X1 inst_cellmath__60_0_I381 (.Y(N679), .A(N508), .B(N513));
NOR2XL inst_cellmath__60_0_I382 (.Y(N680), .A(N514), .B(N517));
NAND2XL inst_cellmath__60_0_I383 (.Y(N681), .A(N514), .B(N517));
NOR2XL inst_cellmath__60_0_I384 (.Y(N682), .A(N518), .B(N521));
NAND2XL inst_cellmath__60_0_I385 (.Y(N683), .A(N518), .B(N521));
NOR2XL inst_cellmath__60_0_I386 (.Y(N684), .A(N523), .B(N522));
NAND2XL inst_cellmath__60_0_I387 (.Y(N685), .A(N523), .B(N522));
NOR2XL inst_cellmath__60_0_I388 (.Y(N686), .A(N525), .B(N524));
NAND2XL inst_cellmath__60_0_I389 (.Y(N687), .A(N525), .B(N524));
NOR2XL inst_cellmath__60_0_I390 (.Y(N688), .A(N414), .B(N526));
NAND2XL inst_cellmath__60_0_I391 (.Y(N689), .A(N414), .B(N526));
AOI21X2 inst_cellmath__60_0_I396 (.Y(N694), .A0(N663), .A1(N660), .B0(N662));
AOI21X2 inst_cellmath__60_0_I400 (.Y(N698), .A0(N667), .A1(N664), .B0(N666));
NAND2X1 inst_cellmath__60_0_I401 (.Y(N699), .A(N667), .B(N665));
AOI21X4 inst_cellmath__60_0_I404 (.Y(N702), .A0(N671), .A1(N668), .B0(N670));
NAND2X4 inst_cellmath__60_0_I405 (.Y(N703), .A(N671), .B(N669));
AOI21X4 inst_cellmath__60_0_I408 (.Y(N706), .A0(N675), .A1(N672), .B0(N674));
NAND2X4 inst_cellmath__60_0_I409 (.Y(N707), .A(N675), .B(N673));
AOI21X1 inst_cellmath__60_0_I412 (.Y(N710), .A0(N679), .A1(N676), .B0(N678));
NAND2X2 inst_cellmath__60_0_I413 (.Y(N711), .A(N679), .B(N677));
AOI21XL inst_cellmath__60_0_I416 (.Y(N714), .A0(N683), .A1(N680), .B0(N682));
NAND2XL inst_cellmath__60_0_I417 (.Y(N715), .A(N683), .B(N681));
INVXL inst_cellmath__60_0_I749 (.Y(N1206), .A(N684));
INVXL inst_cellmath__60_0_I750 (.Y(N1207), .A(N685));
AOI21XL inst_cellmath__60_0_I420 (.Y(N718), .A0(N687), .A1(N684), .B0(N686));
NAND2XL inst_cellmath__60_0_I421 (.Y(N719), .A(N687), .B(N685));
OAI21XL inst_cellmath__60_0_I426 (.Y(N724), .A0(N1207), .A1(N714), .B0(N1206));
OA21X1 inst_cellmath__60_0_I808 (.Y(N1220), .A0(N719), .A1(N714), .B0(N718));
OR2XL inst_cellmath__60_0_I809 (.Y(N1221), .A(N719), .B(N715));
INVX1 inst_cellmath__60_0_I765 (.Y(N1222), .A(N694));
OAI21X2 inst_cellmath__60_0_I444 (.Y(N742), .A0(N699), .A1(N694), .B0(N698));
OAI21X4 inst_cellmath__60_0_I446 (.Y(N744), .A0(N703), .A1(N698), .B0(N702));
NOR2X2 inst_cellmath__60_0_I447 (.Y(N745), .A(N703), .B(N699));
OAI21X2 inst_cellmath__60_0_I448 (.Y(N746), .A0(N707), .A1(N702), .B0(N706));
NOR2XL inst_cellmath__60_0_I449 (.Y(N747), .A(N707), .B(N703));
OAI21X2 inst_cellmath__60_0_I450 (.Y(N748), .A0(N711), .A1(N706), .B0(N710));
NOR2X2 inst_cellmath__60_0_I451 (.Y(N749), .A(N711), .B(N707));
OAI21XL inst_cellmath__60_0_I452 (.Y(N750), .A0(N1221), .A1(N710), .B0(N1220));
NOR2X1 inst_cellmath__60_0_I453 (.Y(N751), .A(N1221), .B(N711));
INVX1 inst_cellmath__60_0_I766 (.Y(N1223), .A(N1222));
INVX1 inst_cellmath__60_0_I767 (.Y(N1224), .A(N742));
AOI21XL inst_cellmath__60_0_I458 (.Y(N756), .A0(N745), .A1(N1222), .B0(N744));
AOI21X1 inst_cellmath__60_0_I460 (.Y(N758), .A0(N747), .A1(N742), .B0(N746));
AOI21X4 inst_cellmath__60_0_I462 (.Y(N760), .A0(N749), .A1(N744), .B0(N748));
NAND2X2 inst_cellmath__60_0_I463 (.Y(N761), .A(N749), .B(N745));
AOI21X2 inst_cellmath__60_0_I464 (.Y(N762), .A0(N751), .A1(N746), .B0(N750));
NAND2XL inst_cellmath__60_0_I465 (.Y(N763), .A(N751), .B(N747));
OAI21X4 inst_cellmath__60_0_I474 (.Y(N772), .A0(N761), .A1(N1223), .B0(N760));
OAI21X2 inst_cellmath__60_0_I476 (.Y(N774), .A0(N763), .A1(N1224), .B0(N762));
INVXL inst_cellmath__60_0_I784 (.Y(N1241), .A(N714));
NAND2BXL inst_cellmath__60_0_I503 (.Y(N801), .AN(N662), .B(N663));
NAND2BXL inst_cellmath__60_0_I506 (.Y(N804), .AN(N664), .B(N665));
NAND2BXL inst_cellmath__60_0_I509 (.Y(N807), .AN(N666), .B(N667));
NAND2BXL inst_cellmath__60_0_I512 (.Y(N810), .AN(N668), .B(N669));
NAND2BXL inst_cellmath__60_0_I515 (.Y(N813), .AN(N670), .B(N671));
NAND2BXL inst_cellmath__60_0_I518 (.Y(N816), .AN(N672), .B(N673));
NAND2BXL inst_cellmath__60_0_I521 (.Y(N819), .AN(N674), .B(N675));
NAND2BXL inst_cellmath__60_0_I524 (.Y(N822), .AN(N676), .B(N677));
NAND2BXL inst_cellmath__60_0_I527 (.Y(N825), .AN(N678), .B(N679));
NAND2BXL inst_cellmath__60_0_I530 (.Y(N828), .AN(N680), .B(N681));
NAND2BXL inst_cellmath__60_0_I533 (.Y(N831), .AN(N682), .B(N683));
NAND2BXL inst_cellmath__60_0_I536 (.Y(N834), .AN(N684), .B(N685));
NAND2BXL inst_cellmath__60_0_I539 (.Y(N837), .AN(N686), .B(N687));
NAND2BXL inst_cellmath__60_0_I542 (.Y(N840), .AN(N688), .B(N689));
NOR2BX1 inst_cellmath__60_0_I838 (.Y(N843), .AN(N1148), .B(N1153));
XOR2XL inst_cellmath__60_0_I811 (.Y(inst_cellmath__60_0_out0[10]), .A(N660), .B(N801));
XNOR2X1 inst_cellmath__60_0_I548 (.Y(inst_cellmath__60_0_out0[11]), .A(N1223), .B(N804));
XNOR2X1 inst_cellmath__60_0_I1545 (.Y(inst_cellmath__60_0_out0[13]), .A(N1224), .B(N810));
XNOR2X1 inst_cellmath__60_0_I813 (.Y(inst_cellmath__60_0_out0[15]), .A(N756), .B(N816));
XNOR2X1 inst_cellmath__60_0_I814 (.Y(inst_cellmath__60_0_out0[17]), .A(N758), .B(N822));
INVXL xor2_A_I868 (.Y(N1253), .A(N772));
MXI2X4 xor2_A_I869 (.Y(inst_cellmath__60_0_out0[19]), .A(N1253), .B(N772), .S0(N828));
XOR2XL inst_cellmath__60_0_I553 (.Y(inst_cellmath__60_0_out0[23]), .A(N774), .B(N840));
XNOR2X1 node_cs_reduced_local_A_I608 (.Y(N852), .A(N807), .B(N665));
XNOR2X1 node_cs_reduced_local_A_I609 (.Y(N853), .A(N807), .B(N664));
MXI2XL inst_cellmath__60_0_I555 (.Y(inst_cellmath__60_0_out0[12]), .A(N852), .B(N853), .S0(N1223));
XNOR2X1 node_cs_reduced_local_A_I610 (.Y(N855), .A(N813), .B(N669));
XNOR2X1 node_cs_reduced_local_A_I611 (.Y(N856), .A(N813), .B(N668));
MXI2XL inst_cellmath__60_0_I557 (.Y(inst_cellmath__60_0_out0[14]), .A(N855), .B(N856), .S0(N1224));
XNOR2X1 node_cs_reduced_local_A_I612 (.Y(N858), .A(N819), .B(N673));
XNOR2X1 node_cs_reduced_local_A_I613 (.Y(N859), .A(N819), .B(N672));
MXI2XL inst_cellmath__60_0_I559 (.Y(inst_cellmath__60_0_out0[16]), .A(N858), .B(N859), .S0(N756));
XNOR2X1 node_cs_reduced_local_A_I614 (.Y(N861), .A(N825), .B(N677));
XNOR2X1 node_cs_reduced_local_A_I615 (.Y(N862), .A(N825), .B(N676));
MXI2XL inst_cellmath__60_0_I561 (.Y(inst_cellmath__60_0_out0[18]), .A(N861), .B(N862), .S0(N758));
XNOR2X1 node_cs_reduced_local_A_I616 (.Y(N864), .A(N831), .B(N681));
XNOR2X1 node_cs_reduced_local_A_I617 (.Y(N865), .A(N831), .B(N680));
MXI2XL inst_cellmath__60_0_I563 (.Y(inst_cellmath__60_0_out0[20]), .A(N865), .B(N864), .S0(N772));
XNOR2X1 node_cs_local_A_I618 (.Y(N867), .A(N834), .B(N1241));
NOR2BX1 node_cs_local_A_I815 (.Y(N1057), .AN(N715), .B(N1241));
XOR2XL node_cs_local_A_I620 (.Y(N868), .A(N834), .B(N1057));
MXI2XL inst_cellmath__60_0_I565 (.Y(inst_cellmath__60_0_out0[21]), .A(N867), .B(N868), .S0(N772));
XNOR2X1 node_cs_local_A_I621 (.Y(N870), .A(N837), .B(N724));
NOR2XL andori2bb1_A_I870 (.Y(N1260), .A(N1207), .B(N715));
NOR2XL andori2bb1_A_I871 (.Y(N1066), .A(N1260), .B(N724));
XOR2XL node_cs_local_A_I623 (.Y(N871), .A(N837), .B(N1066));
MXI2XL inst_cellmath__60_0_I567 (.Y(inst_cellmath__60_0_out0[22]), .A(N870), .B(N871), .S0(N772));
XNOR2X1 node_cs_reduced_local_A_I624 (.Y(N873), .A(N843), .B(N689));
XNOR2X1 node_cs_reduced_local_A_I625 (.Y(N874), .A(N843), .B(N688));
MXI2XL inst_cellmath__60_0_I569 (.Y(inst_cellmath__60_0_out0[24]), .A(N874), .B(N873), .S0(N774));
assign inst_cellmath__60_0_out0[1] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_noninc_a_cellmath__55_2WWMM_bdw1471647203_bdw (
	inst_noninc_a_cellmath__55_2WWMM_out0,
	inst_noninc_a_cellmath__55_2WWMM_in0
	); /* architecture "gate_level" */ 
output [52:0] inst_noninc_a_cellmath__55_2WWMM_out0;
input [22:16] inst_noninc_a_cellmath__55_2WWMM_in0;
wire N1044,N1045,N1060,N1061,N1062,N1066,N1068 
	,N1084,N1086,N1089,N1092,N1093,N1102,N1103,N2138 
	,N2140,N2141,N2142,N2146,N2147,N2163,N2166,N2168 
	,N2170,N2174,N2175,N2176,N2179,N2180,N2199,N2200 
	,N2201,N2202,N2203,N2211,N2212,N2213,N2214,N2215 
	,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223 
	,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243 
	,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251 
	,N2253,N2256,N2257,N2258,N2259,N2261,N3281,N3282 
	,N3287,N3304,N3305,N3306,N3309,N3314,N3322,N3327 
	,N4329,N4342,N4344,N4345,N4346,N4350,N4351,N4367 
	,N4371,N4376,N4377,N4380,N4382,N4396,N4411,N4413 
	,N4414,N4415,N4416,N4417,N4425,N4426,N4427,N4428 
	,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436 
	,N4437,N4448,N4449,N4450,N4451,N4452,N4453,N4454 
	,N4455,N4456,N4457,N4458,N4459,N4461,N4462,N4463 
	,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4473 
	,N4478,N4479,N4480,N4481,N4482,N4483,N4493,N4494 
	,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502 
	,N4503,N4504,N4505,N4506,N4507,N4513,N4514,N4515 
	,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523 
	,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531 
	,N4532,N4533,N4534,N4535,N5537,N5550,N5553,N5554 
	,N5555,N5558,N5578,N5584,N5586,N5591,N5592,N5593 
	,N5594,N6610,N6613,N6633,N6635,N6638,N6641,N6642 
	,N6643,N6648,N6657,N6670,N6671,N6672,N6673,N6683 
	,N6684,N6685,N6686,N6687,N6690,N6691,N6692,N6693 
	,N6694,N6695,N6696,N6697,N6698,N6707,N6708,N6709 
	,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717 
	,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725 
	,N6726,N6727,N7736,N7739,N7753,N7755,N7759,N7780 
	,N7783,N7790,N7795,N7799,N8814,N8819,N8831,N8843 
	,N8845,N8861,N8862,N8863,N8867,N8868,N8870,N8871 
	,N8873,N8895,N8896,N8897,N8898,N8899,N8900,N8901 
	,N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916 
	,N8917,N8919,N8922,N8923,N8924,N8925,N8926,N8933 
	,N8934,N8935,N8936,N8937,N8938,N8939,N8940,N8941 
	,N8942,N8943,N8944,N8945,N8946,N8947,N8948,N8949 
	,N8950,N8951,N8952,N8953,N8954,N8962,N8963,N8964 
	,N8965,N8966,N8967,N8968,N8972,N8977,N8978,N8979 
	,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987 
	,N8988,N8989,N8990,N8991,N8998,N8999,N9000,N9001 
	,N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009 
	,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017 
	,N9018,N9019,N9020,N9022,N9028,N9029,N9030,N9031 
	,N9032,N9033,N9034,N9036,N9039,N9042,N9043,N9044 
	,N9045,N9046,N9047,N9048,N9049,N9050,N9051,N9052 
	,N9053,N9054,N9055,N9056,N9057,N9063,N9064,N9065 
	,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073 
	,N9074,N9075,N9076,N9077,N9078,N9079,N9080,N9081 
	,N9082,N9083,N9084,N9085,N9086,N10112,N10134,N10137 
	,N10146,N11159,N11176,N11178,N11181,N11204,N11207,N11210 
	,N11236,N11237,N11238,N11239,N11240,N11241,N11242,N11243 
	,N11248,N11249,N11250,N11251,N11252,N11253,N11254,N11255 
	,N11256,N11257,N11258,N11259,N11271,N11272,N11273,N11274 
	,N11275,N11276,N11277,N11278,N11279,N11280,N11281,N11282 
	,N11283,N11284,N11285,N11286,N11287,N11292,N11293,N11294 
	,N11295,N11296,N12316,N12319,N12328,N12343,N12346,N12357 
	,N12362,N12363,N12366,N12367,N13404,N13406,N13407,N13408 
	,N13411,N13437,N13443,N13448,N13459,N13462,N13471,N13472 
	,N13473,N13477,N13478,N13487,N13488,N13489,N13490,N13491 
	,N13492,N13493,N13494,N13495,N13496,N13497,N13498,N13499 
	,N13501,N13508,N13509,N13510,N13511,N13512,N13513,N13514 
	,N13515,N13516,N13517,N13518,N13519,N13520,N13521,N13522 
	,N13523,N13524,N13525,N13526,N13527,N13528,N13529,N13538 
	,N13539,N13540,N13541,N13542,N13543,N13544,N13545,N13546 
	,N13551,N13552,N13553,N13554,N13555,N13556,N13557,N13558 
	,N13559,N13560,N13561,N13562,N13563,N13564,N13565,N13566 
	,N13567,N13569,N13572,N13573,N13574,N13575,N13576,N13577 
	,N13578,N13579,N13580,N13581,N13582,N13583,N13584,N13585 
	,N13586,N13587,N13588,N13589,N13590,N13591,N13592,N13593 
	,N13594,N14617,N14619,N14621,N14638,N14641,N14649,N14658 
	,N15695,N15708,N15724,N15725,N15750,N15751,N15752,N15753 
	,N15754,N15755,N15756,N15762,N15763,N15764,N15765,N15766 
	,N15767,N15768,N15769,N15770,N15771,N15772,N15773,N15774 
	,N15775,N15776,N15783,N15784,N15785,N15786,N15787,N15788 
	,N15789,N15790,N15791,N15792,N15793,N15794,N15795,N15796 
	,N15797,N15798,N15799,N15800,N15801,N15802,N15804,N15805 
	,N16832,N16845,N16861,N16862,N16869,N16878,N16879,N16882 
	,N17901,N17908,N17948,N17951,N17969,N17970,N17971,N17972 
	,N17973,N17974,N17975,N17976,N17982,N17983,N17984,N17985 
	,N17986,N17987,N17989,N17990,N17991,N17992,N17993,N17994 
	,N17995,N17996,N17997,N17998,N18002,N18003,N18004,N18005 
	,N18006,N18007,N18008,N18009,N18010,N18011,N18012,N18013 
	,N18014,N18015,N18016,N18017,N18018,N18019,N18020,N18023 
	,N18024,N18025,N18026,N18034,N18035,N18036,N18037,N18038 
	,N18039,N18040,N18041,N18046,N18047,N18048,N18049,N18050 
	,N18051,N18052,N18053,N18054,N18055,N18056,N18057,N18058 
	,N18059,N18060,N18061,N18062,N18067,N18068,N18069,N18070 
	,N18071,N18072,N18073,N18074,N18075,N18076,N18077,N18078 
	,N18079,N18080,N18081,N18082,N18083,N18084,N18085,N18086 
	,N18087,N18088,N18089,N18090,N18094,N18095,N18096,N18097 
	,N18098,N18099,N18100,N18101,N18102,N18103,N18106,N18107 
	,N18108,N18109,N18110,N18111,N18112,N18113,N18114,N18115 
	,N18116,N18117,N18118,N18119,N18120,N18121,N18122,N18125 
	,N18126,N18127,N18128,N18129,N18130,N18131,N18132,N18133 
	,N18134,N18135,N18136,N18137,N18138,N18139,N18140,N18141 
	,N18142,N18143,N18144,N18145,N18146,N18147,N18148,N18213 
	,N18215,N18217,N18219,N18221,N18229,N18231,N18233,N18235 
	,N18239,N18241,N18243,N18245,N18247,N18249,N18251,N18253 
	,N18259,N18261,N18265,N18269,N18273,N18275,N18277,N18279 
	,N18281,N18283,N18287,N18289,N18291,N18293,N18295,N18297 
	,N18301,N18307,N18309,N18311,N18315,N18319,N18321,N18323 
	,N18327,N18329,N18331,N18333,N18335,N18337,N18339,N18341 
	,N18343,N18347,N18349,N18351,N18353,N18357,N18359,N18361 
	,N18397,N18398,N18399,N18400,N18403,N18405,N18406,N18407 
	,N18409,N18410,N18411,N18415,N18418,N18420,N18430,N18432 
	,N18435,N18439,N18440,N18445,N18448,N18450,N18454,N18455 
	,N18458,N18460,N18465,N18466,N18467,N18470,N18474,N18476 
	,N18477,N18478,N18479,N18483,N18489,N18495,N18496,N18498 
	,N18501,N18508,N18510,N18514,N18531,N18545,N18546,N18547 
	,N18569,N18570,N18572,N18573,N18578,N18579,N18580,N18583 
	,N18596,N18601,N18608,N18609,N18610,N18672,N18677,N18702 
	,N18705,N18706,N18707,N18717,N18722,N18725,N18728,N18729 
	,N18730,N18735,N18739,N18747,N18748,N18802,N18820,N18831 
	,N18832,N18833,N18834,N18865,N18880,N18884,N18885,N18889 
	,N18890,N18892,N18893,N18896,N18897,N18901,N18902,N18905 
	,N18906,N18907,N18908,N18909,N18911,N18931,N18933,N18937 
	,N18950,N18953,N19038,N19085,N19086,N19107,N19111,N19112 
	,N19132,N19139,N19146,N19153,N19160,N21286;
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14213 (.Y(N18884), .A(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I14214 (.Y(N18885), .A(N18884));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13729 (.Y(N18400), .A(N18885));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13728 (.Y(N18399), .A(N18885));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13727 (.Y(N18398), .A(N18885));
CLKINVX8 inst_noninc_a_cellmath__55_2WWMM_I13726 (.Y(N18397), .A(N18885));
CLKINVX8 inst_noninc_a_cellmath__55_2WWMM_I14225 (.Y(N18896), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I14226 (.Y(N18897), .A(N18896));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I13735 (.Y(N18406), .A(N18897));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13734 (.Y(N18405), .A(N18897));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13732 (.Y(N18403), .A(N18897));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14219 (.Y(N18890), .A(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I14222 (.Y(N18893), .A(N18890));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I322 (.Y(N18213), .A0(N18893), .A1(N18406), .B0(N18397), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13736 (.Y(N18407), .A(N18213));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13740 (.Y(N18411), .A(N18407));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13739 (.Y(N18410), .A(N18407));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13738 (.Y(N18409), .A(N18407));
NAND2X4 inst_noninc_a_cellmath__55_2WWMM_I323 (.Y(N18215), .A(N18406), .B(N18397));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13744 (.Y(N18415), .A(N18215));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I13749 (.Y(N18420), .A(N18415));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13747 (.Y(N18418), .A(N18415));
NAND2X2 inst_noninc_a_cellmath__55_2WWMM_I333 (.Y(N18217), .A(N18406), .B(N18893));
INVXL buf1_A_I16716 (.Y(N21286), .A(N18217));
INVXL buf1_A_I16717 (.Y(N18432), .A(N21286));
BUFX6 inst_noninc_a_cellmath__55_2WWMM_I16699 (.Y(N18430), .A(N18217));
NOR2X2 inst_noninc_a_cellmath__55_2WWMM_I334 (.Y(N18219), .A(N18406), .B(N18397));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13764 (.Y(N18435), .A(N18219));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13769 (.Y(N18440), .A(N18435));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13768 (.Y(N18439), .A(N18435));
NAND2X2 inst_noninc_a_cellmath__55_2WWMM_I339 (.Y(N18221), .A(N18893), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13774 (.Y(N18445), .A(N18221));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13779 (.Y(N18450), .A(N18445));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13777 (.Y(N18448), .A(N18445));
NOR2X2 inst_noninc_a_cellmath__55_2WWMM_I14567 (.Y(N18454), .A(N18403), .B(N18893));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13784 (.Y(N18455), .A(N18454));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13789 (.Y(N18460), .A(N18455));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13787 (.Y(N18458), .A(N18455));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14221 (.Y(N18892), .A(N18890));
OR2X1 inst_noninc_a_cellmath__55_2WWMM_I14477 (.Y(N18465), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B(N18892));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13799 (.Y(N18470), .A(N18465));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13796 (.Y(N18467), .A(N18465));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13795 (.Y(N18466), .A(N18465));
OR2X6 inst_noninc_a_cellmath__55_2WWMM_I14478 (.Y(N18474), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B(N18397));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13808 (.Y(N18479), .A(N18474));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13807 (.Y(N18478), .A(N18474));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13806 (.Y(N18477), .A(N18474));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13805 (.Y(N18476), .A(N18474));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14234 (.Y(N18905), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14235 (.Y(N18906), .A(N18905));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I14236 (.Y(N18907), .A(N18906));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I14237 (.Y(N18908), .A(N18907));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I13812 (.Y(N18483), .A(N18908));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I13837 (.Y(N18508), .A(N18483));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I13825 (.Y(N18496), .A(N18483));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I13860 (.Y(N18531), .A(N18908));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13843 (.Y(N18514), .A(N18508));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I13839 (.Y(N18510), .A(N18508));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13830 (.Y(N18501), .A(N18496));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13827 (.Y(N18498), .A(N18496));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13824 (.Y(N18495), .A(N18496));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13818 (.Y(N18489), .A(N18508));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14231 (.Y(N18902), .A(N18896));
BUFX2 inst_noninc_a_cellmath__55_2WWMM_I14526 (.Y(N18950), .A(N18905));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I14282 (.Y(N18953), .A(N18950));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I749 (.Y(N18229), .A0(N18531), .A1(N18215), .B0(N18902), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I750 (.Y(N1044), .A0(N18531), .A1(N18454), .B0(N18410), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I751 (.Y(N1045), .A0(N18531), .A1(N18448), .B0(N18215), .B1(N18953));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I752 (.Y(N18231), .A(N18953), .B(N18219));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I759 (.Y(N1060), .A0(N18531), .A1(N18219), .B0(N18902), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I760 (.Y(N1061), .A0(N18531), .A1(N18403), .B0(N18892), .B1(N18953));
INVXL inst_noninc_a_cellmath__55_2WWMM_I761 (.Y(N1062), .A(N18430));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I762 (.Y(N18233), .A0(N18531), .A1(N18432), .B0(N18219), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I763 (.Y(N18235), .A0(N18531), .A1(N18902), .B0(N18892), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I765 (.Y(N1066), .A0(N18531), .A1(N18454), .B0(N18440), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I766 (.Y(N18239), .A0(N18531), .A1(N18403), .B0(N18440), .B1(N18953));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13874 (.Y(N18545), .A(N18239));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13876 (.Y(N18547), .A(N18545));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13875 (.Y(N18546), .A(N18545));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I767 (.Y(N1068), .A(N18531), .B(N18221));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I777 (.Y(N1084), .A0(N18531), .A1(N18454), .B0(N18430), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I779 (.Y(N1086), .A0(N18531), .A1(N18892), .B0(N18440), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I780 (.Y(N18241), .A0(N18531), .A1(N18448), .B0(N18430), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I781 (.Y(N18243), .A0(N18531), .A1(N18470), .B0(N18902), .B1(N18953));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I782 (.Y(N1089), .A(N18953), .B(N18460));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I783 (.Y(N1092), .A0(N18531), .A1(N18892), .B0(N18418), .B1(N18953));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I784 (.Y(N1093), .A(N18531), .B(N18219));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I785 (.Y(N18245), .A(N18953), .B(N18479));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I786 (.Y(N18247), .A(N18953), .B(N18902));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I788 (.Y(N1102), .A0(N18531), .A1(N18403), .B0(N18902), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I789 (.Y(N1103), .A0(N18531), .A1(N18219), .B0(N18418), .B1(N18953));
NAND2X4 inst_noninc_a_cellmath__55_2WWMM_I1133 (.Y(N18249), .A(N18397), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I1136 (.Y(N18251), .A0(N18403), .A1(N18397), .B0(N18893), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13898 (.Y(N18569), .A(N18251));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I13902 (.Y(N18573), .A(N18569));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13901 (.Y(N18572), .A(N18569));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I13899 (.Y(N18570), .A(N18569));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I1551 (.Y(N18253), .A(N18489), .B(N18466));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14230 (.Y(N18901), .A(N18896));
AO22XL inst_noninc_a_cellmath__55_2WWMM_I14554 (.Y(N18578), .A0(N18403), .A1(N18953), .B0(N18489), .B1(N18901));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13909 (.Y(N18580), .A(N18578));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13908 (.Y(N18579), .A(N18578));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I14485 (.Y(N18583), .A(N18901), .B(N18953));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I1561 (.Y(N18259), .A0(N18489), .A1(N18570), .B0(N18249), .B1(N18953));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1562 (.Y(N2138), .A(N18489), .B(N18397));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1563 (.Y(N2140), .A0(N18489), .A1(N18410), .B0(N18448), .B1(N18953));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1564 (.Y(N2141), .A0(N18448), .A1(N18489), .B0(N18570), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1565 (.Y(N2142), .A0(N18489), .A1(N18440), .B0(N18570), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1566 (.Y(N18261), .A0(N18489), .A1(N18893), .B0(N18410), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1569 (.Y(N2146), .A0(N18489), .A1(N18570), .B0(N18440), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1570 (.Y(N2147), .A0(N18510), .A1(N18249), .B0(N18478), .B1(N18953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1572 (.Y(N18265), .A0(N18510), .A1(N18420), .B0(N18466), .B1(N18953));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I14491 (.Y(N18596), .A(N18953), .B(N18420));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1574 (.Y(N18269), .A(N18510), .B(N18467));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1580 (.Y(N2163), .A(N18397), .B(N18953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I14556 (.Y(N18601), .A0(N18466), .A1(N18953), .B0(N18510), .B1(N18901));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1582 (.Y(N2166), .A0(N18510), .A1(N18467), .B0(N18432), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1583 (.Y(N18273), .A0(N18901), .A1(N18489), .B0(N18478), .B1(N18953));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1584 (.Y(N2168), .A(N18489), .B(N18901));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1585 (.Y(N2170), .A(N18489), .B(N18893));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1588 (.Y(N2174), .A0(N18489), .A1(N18420), .B0(N18249), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1589 (.Y(N2175), .A0(N18901), .A1(N18489), .B0(N18460), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1590 (.Y(N2176), .A0(N18489), .A1(N18460), .B0(N18249), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1592 (.Y(N18275), .A0(N18902), .A1(N18489), .B0(N18410), .B1(N18953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1593 (.Y(N2179), .A0(N18489), .A1(N18570), .B0(N18432), .B1(N18953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1594 (.Y(N2180), .A0(N18489), .A1(N18440), .B0(N18466), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1596 (.Y(N18277), .A0(N18489), .A1(N18397), .B0(N18249), .B1(N18953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1597 (.Y(N18279), .A0(N18498), .A1(N18410), .B0(N18430), .B1(N18953));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13937 (.Y(N18608), .A(N18279));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13939 (.Y(N18610), .A(N18608));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13938 (.Y(N18609), .A(N18608));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1598 (.Y(N18281), .A0(N18467), .A1(N18498), .B0(N18215), .B1(N18953));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I14001 (.Y(N18672), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14006 (.Y(N18677), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1605 (.Y(N2199), .A0(N18672), .A1(N18253), .B0(N18229), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1606 (.Y(N2200), .A0(N18672), .A1(N18398), .B0(N1044), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1607 (.Y(N2201), .A0(N18672), .A1(N18902), .B0(N1045), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1608 (.Y(N2202), .A0(N18672), .A1(N18580), .B0(N18231), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1609 (.Y(N2203), .A(N18672), .B(N18583));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1615 (.Y(N2211), .A0(N18672), .A1(N18259), .B0(N1060), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1616 (.Y(N2212), .A0(N18672), .A1(N2138), .B0(N1061), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1617 (.Y(N2213), .A0(N18672), .A1(N2140), .B0(N1062), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1618 (.Y(N2214), .A0(N18672), .A1(N2141), .B0(N18233), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1619 (.Y(N2215), .A0(N18672), .A1(N2142), .B0(N18235), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1620 (.Y(N2216), .A0(N18672), .A1(N18261), .B0(N18407), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1621 (.Y(N2217), .A0(N18672), .A1(N18235), .B0(N1066), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1622 (.Y(N2218), .A0(N18672), .A1(N18261), .B0(N18547), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1623 (.Y(N2219), .A0(N18672), .A1(N2146), .B0(N1068), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1624 (.Y(N2220), .A0(N18672), .A1(N2147), .B0(N18893), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1625 (.Y(N2221), .A0(N18672), .A1(N18569), .B0(N18902), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14238 (.Y(N18909), .A(N18907));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1626 (.Y(N2222), .A0(N18672), .A1(N18265), .B0(N18909), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1627 (.Y(N2223), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18596));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1628 (.Y(N18283), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18269));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1633 (.Y(N2236), .A0(N18672), .A1(N18247), .B0(N1084), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1634 (.Y(N2237), .A0(N18672), .A1(N2163), .B0(N18233), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1635 (.Y(N2238), .A0(N18672), .A1(N18601), .B0(N1086), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1636 (.Y(N2239), .A0(N18672), .A1(N2166), .B0(N18241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1637 (.Y(N2240), .A0(N18672), .A1(N18273), .B0(N18243), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1638 (.Y(N2241), .A0(N18672), .A1(N2168), .B0(N1089), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1639 (.Y(N2242), .A0(N18672), .A1(N2170), .B0(N1092), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1640 (.Y(N2243), .A0(N18672), .A1(N18243), .B0(N1093), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1641 (.Y(N2244), .A0(N18672), .A1(N18601), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1642 (.Y(N2245), .A0(N18672), .A1(N2174), .B0(N18247), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1643 (.Y(N2246), .A0(N18672), .A1(N2175), .B0(N18407), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1644 (.Y(N2247), .A0(N18672), .A1(N2176), .B0(N1102), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1645 (.Y(N2248), .A0(N18672), .A1(N18273), .B0(N1103), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1646 (.Y(N2249), .A0(N18672), .A1(N18275), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1647 (.Y(N2250), .A0(N18672), .A1(N2179), .B0(N18247), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1648 (.Y(N2251), .A(N18672), .B(N2180));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1649 (.Y(N2253), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1650 (.Y(N2256), .A0(N18672), .A1(N18277), .B0(N18397), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1651 (.Y(N2257), .A0(N18672), .A1(N18610), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1652 (.Y(N2258), .A0(N18672), .A1(N18281), .B0(N18489), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1653 (.Y(N2259), .A(N18672), .B(N18269));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1654 (.Y(N2261), .A(N18672), .B(N18596));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I14497 (.Y(N18702), .A(N18498), .B(N18403));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2417 (.Y(N18287), .A0(N18498), .A1(N18420), .B0(N18460), .B1(N18953));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I2418 (.Y(N18289), .A0(N18498), .A1(N18460), .B0(N18478), .B1(N18953));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14034 (.Y(N18705), .A(N18289));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14036 (.Y(N18707), .A(N18705));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14035 (.Y(N18706), .A(N18705));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2419 (.Y(N3281), .A0(N18495), .A1(N18448), .B0(N18249), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2420 (.Y(N3282), .A0(N18495), .A1(N18467), .B0(N18893), .B1(N18953));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2423 (.Y(N3287), .A(N18953), .B(N18470));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14218 (.Y(N18889), .A(N18884));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I2424 (.Y(N18291), .A0(N18495), .A1(N18889), .B0(N18398), .B1(N18953));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I2425 (.Y(N18293), .A0(N18495), .A1(N18573), .B0(N18403), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2426 (.Y(N18295), .A0(N18495), .A1(N18249), .B0(N18398), .B1(N18953));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I2427 (.Y(N18297), .A0(N18501), .A1(N18409), .B0(N18902), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I14500 (.Y(N18717), .A0(N18403), .A1(N18953), .B0(N18501), .B1(N18440));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I2429 (.Y(N18301), .A(N18501), .B(N18448));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2435 (.Y(N3304), .A0(N18501), .A1(N18889), .B0(N18467), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2436 (.Y(N3305), .A0(N18501), .A1(N18478), .B0(N18448), .B1(N18953));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2437 (.Y(N3306), .A(N18495), .B(N18420));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2438 (.Y(N3309), .A(N18953), .B(N18448));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I14502 (.Y(N18722), .A0(N18889), .A1(N18953), .B0(N18495), .B1(N18573));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2441 (.Y(N3314), .A0(N18249), .A1(N18495), .B0(N18410), .B1(N18953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I14504 (.Y(N18725), .A0(N18953), .A1(N18570), .B0(N18430), .B1(N18495));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2448 (.Y(N3322), .A0(N18495), .A1(N18249), .B0(N18902), .B1(N18953));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14260 (.Y(N18931), .A(N18906));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14266 (.Y(N18937), .A(N18931));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I2449 (.Y(N18307), .A0(N18495), .A1(N18440), .B0(N18398), .B1(N18937));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I2450 (.Y(N18309), .A0(N18495), .A1(N18476), .B0(N18409), .B1(N18937));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14057 (.Y(N18728), .A(N18309));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14059 (.Y(N18730), .A(N18728));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14058 (.Y(N18729), .A(N18728));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2452 (.Y(N18311), .A0(N18495), .A1(N18889), .B0(N18460), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2453 (.Y(N3327), .A0(N18403), .A1(N18495), .B0(N18409), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I14561 (.Y(N18735), .A0(N18420), .A1(N18937), .B0(N18495), .B1(N18405));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3210 (.Y(N4329), .A0(N18498), .A1(N18398), .B0(N18889), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I3219 (.Y(N4342), .A0(N18498), .A1(N18439), .B0(N18448), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3220 (.Y(N18315), .A0(N18498), .A1(N18420), .B0(N18405), .B1(N18937));
INVXL inst_noninc_a_cellmath__55_2WWMM_I3221 (.Y(N4344), .A(N18418));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3222 (.Y(N4345), .A0(N18498), .A1(N18476), .B0(N18439), .B1(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3223 (.Y(N4346), .A(N18470), .B(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I14509 (.Y(N18739), .A(N18498), .B(N18249));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3225 (.Y(N4350), .A0(N18498), .A1(N18405), .B0(N18398), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I3226 (.Y(N4351), .A0(N18498), .A1(N18405), .B0(N18573), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I3228 (.Y(N18319), .A0(N18498), .A1(N18460), .B0(N18573), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3229 (.Y(N18321), .A0(N18498), .A1(N18430), .B0(N18476), .B1(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3231 (.Y(N18323), .A(N18420), .B(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3237 (.Y(N4367), .A(N18498), .B(N18889));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3239 (.Y(N4371), .A(N18501), .B(N18430));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3241 (.Y(N4376), .A0(N18501), .A1(N18889), .B0(N18249), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I3242 (.Y(N4377), .A0(N18501), .A1(N18439), .B0(N18430), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3245 (.Y(N4380), .A0(N18501), .A1(N18249), .B0(N18448), .B1(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3247 (.Y(N4382), .A(N18501), .B(N18476));
AO22XL inst_noninc_a_cellmath__55_2WWMM_I16706 (.Y(N18747), .A0(N18460), .A1(N18937), .B0(N18501), .B1(N18249));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14077 (.Y(N18748), .A(N18747));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3255 (.Y(N4396), .A0(N18902), .A1(N18501), .B0(N18573), .B1(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3256 (.Y(N18327), .A(N18501), .B(N18439));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3263 (.Y(N4411), .A(N18677), .B(N2168));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3264 (.Y(N4413), .A0(N18677), .A1(N4329), .B0(N18398), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3265 (.Y(N4414), .A0(N18677), .A1(N18293), .B0(N18901), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3266 (.Y(N4415), .A0(N18677), .A1(N18717), .B0(N18579), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3267 (.Y(N4416), .A0(N18677), .A1(N18583), .B0(N18702), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3268 (.Y(N4417), .A(N18672), .B(N18583));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3273 (.Y(N4425), .A0(N18672), .A1(N4342), .B0(N18287), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3274 (.Y(N4426), .A0(N18672), .A1(N18315), .B0(N18707), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3275 (.Y(N4427), .A0(N18672), .A1(N4344), .B0(N3281), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3276 (.Y(N4428), .A0(N18672), .A1(N4345), .B0(N3282), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3277 (.Y(N4429), .A0(N18672), .A1(N4346), .B0(N18241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3278 (.Y(N4430), .A0(N18672), .A1(N18739), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3279 (.Y(N4431), .A0(N18672), .A1(N4350), .B0(N3287), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3280 (.Y(N4432), .A0(N18672), .A1(N4351), .B0(N18291), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3281 (.Y(N4433), .A0(N18672), .A1(N2179), .B0(N18293), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3282 (.Y(N4434), .A0(N18672), .A1(N18319), .B0(N18295), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3283 (.Y(N4435), .A0(N18672), .A1(N18321), .B0(N18297), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3284 (.Y(N4436), .A0(N18672), .A1(N18735), .B0(N18717), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3285 (.Y(N4437), .A0(N18672), .A1(N18323), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3286 (.Y(N18329), .A(N18672), .B(N18323));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3291 (.Y(N4448), .A0(N18672), .A1(N4367), .B0(N3304), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3292 (.Y(N4449), .A0(N18672), .A1(N18722), .B0(N3305), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3293 (.Y(N4450), .A0(N18672), .A1(N4371), .B0(N3306), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3294 (.Y(N4451), .A0(N18672), .A1(N18253), .B0(N3309), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3295 (.Y(N4452), .A0(N18672), .A1(N4376), .B0(N18233), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3296 (.Y(N4453), .A0(N18672), .A1(N4377), .B0(N18722), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3297 (.Y(N4454), .A0(N18672), .A1(N2174), .B0(N3314), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3298 (.Y(N4455), .A0(N18672), .A1(N18287), .B0(N18241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3299 (.Y(N4456), .A0(N18672), .A1(N4380), .B0(N18546), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3300 (.Y(N4457), .A0(N18672), .A1(N18311), .B0(N18725), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3301 (.Y(N4458), .A0(N18677), .A1(N4382), .B0(N18725), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2BXL inst_noninc_a_cellmath__55_2WWMM_I14511 (.Y(N4459), .AN(N18747), .B(N18677));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3303 (.Y(N4461), .A0(N18677), .A1(N18229), .B0(N3282), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3304 (.Y(N4462), .A0(N18677), .A1(N18901), .B0(N3322), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3305 (.Y(N4463), .A0(N18247), .A1(N18677), .B0(N18307), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3306 (.Y(N4464), .A0(N18677), .A1(N18398), .B0(N18730), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3307 (.Y(N4465), .A0(N18677), .A1(N18405), .B0(N18601), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3308 (.Y(N4466), .A0(N18677), .A1(N18291), .B0(N18311), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3309 (.Y(N4467), .A0(N18677), .A1(N4396), .B0(N3327), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3310 (.Y(N4468), .A0(N18677), .A1(N18327), .B0(N18735), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3311 (.Y(N4469), .A0(N18677), .A1(N18909), .B0(N18247), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3312 (.Y(N4470), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18908));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3313 (.Y(N4473), .A(N18677), .B(N18501));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14367 (.Y(N19038), .A(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14415 (.Y(N19086), .A(N19038));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I14131 (.Y(N18802), .A(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3317 (.Y(N4478), .A0(N18802), .A1(N4411), .B0(N2199), .B1(N19086));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14414 (.Y(N19085), .A(N19038));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3318 (.Y(N4479), .A0(N18802), .A1(N4413), .B0(N2200), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3319 (.Y(N4480), .A0(N18802), .A1(N4414), .B0(N2201), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3320 (.Y(N4481), .A0(N18802), .A1(N4415), .B0(N2202), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3321 (.Y(N4482), .A0(N18802), .A1(N4416), .B0(N2203), .B1(N19085));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3322 (.Y(N4483), .A(N19085), .B(N4417));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3327 (.Y(N4493), .A0(N18802), .A1(N4425), .B0(N2211), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3328 (.Y(N4494), .A0(N18802), .A1(N4426), .B0(N2212), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3329 (.Y(N4495), .A0(N18802), .A1(N4427), .B0(N2213), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3330 (.Y(N4496), .A0(N18802), .A1(N4428), .B0(N2214), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3331 (.Y(N4497), .A0(N18802), .A1(N4429), .B0(N2215), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3332 (.Y(N4498), .A0(N18802), .A1(N4430), .B0(N2216), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3333 (.Y(N4499), .A0(N18802), .A1(N4431), .B0(N2217), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3334 (.Y(N4500), .A0(N18802), .A1(N4432), .B0(N2218), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3335 (.Y(N4501), .A0(N18802), .A1(N4433), .B0(N2219), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3336 (.Y(N4502), .A0(N18802), .A1(N4434), .B0(N2220), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3337 (.Y(N4503), .A0(N18802), .A1(N4435), .B0(N2221), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3338 (.Y(N4504), .A0(N18802), .A1(N4436), .B0(N2222), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3339 (.Y(N4505), .A0(N18802), .A1(N4437), .B0(N2223), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3340 (.Y(N4506), .A0(N18802), .A1(N18329), .B0(N18283), .B1(N19085));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3341 (.Y(N4507), .A(N18802), .B(N2253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3345 (.Y(N4513), .A0(N18802), .A1(N4448), .B0(N2236), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3346 (.Y(N4514), .A0(N18802), .A1(N4449), .B0(N2237), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3347 (.Y(N4515), .A0(N18802), .A1(N4450), .B0(N2238), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3348 (.Y(N4516), .A0(N18802), .A1(N4451), .B0(N2239), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3349 (.Y(N4517), .A0(N18802), .A1(N4452), .B0(N2240), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3350 (.Y(N4518), .A0(N18802), .A1(N4453), .B0(N2241), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3351 (.Y(N4519), .A0(N18802), .A1(N4454), .B0(N2242), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3352 (.Y(N4520), .A0(N18802), .A1(N4455), .B0(N2243), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3353 (.Y(N4521), .A0(N18802), .A1(N4456), .B0(N2244), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3354 (.Y(N4522), .A0(N18802), .A1(N4457), .B0(N2245), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3355 (.Y(N4523), .A0(N18802), .A1(N4458), .B0(N2246), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3356 (.Y(N4524), .A0(N18802), .A1(N4459), .B0(N2247), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3357 (.Y(N4525), .A0(N18802), .A1(N4461), .B0(N2248), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3358 (.Y(N4526), .A0(N18802), .A1(N4462), .B0(N2249), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3359 (.Y(N4527), .A0(N18802), .A1(N4463), .B0(N2250), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3360 (.Y(N4528), .A0(N18802), .A1(N4464), .B0(N2251), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3361 (.Y(N4529), .A0(N18802), .A1(N4465), .B0(N2253), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3362 (.Y(N4530), .A0(N18802), .A1(N4466), .B0(N2256), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3363 (.Y(N4531), .A0(N18802), .A1(N4467), .B0(N2257), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3364 (.Y(N4532), .A0(N18802), .A1(N4468), .B0(N2258), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3365 (.Y(N4533), .A0(N18802), .A1(N4469), .B0(N2259), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3366 (.Y(N4534), .A0(N18802), .A1(N4470), .B0(N2261), .B1(N19085));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3367 (.Y(N4535), .A(N19085), .B(N4473));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I14262 (.Y(N18933), .A(N18931));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4119 (.Y(N18331), .A0(N18501), .A1(N18477), .B0(N18430), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4121 (.Y(N5537), .A0(N18501), .A1(N18249), .B0(N18430), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4129 (.Y(N5550), .A0(N18501), .A1(N18439), .B0(N18460), .B1(N18933));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4131 (.Y(N18333), .A0(N18501), .A1(N18249), .B0(N18889), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4132 (.Y(N5553), .A0(N18501), .A1(N18398), .B0(N18439), .B1(N18933));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4133 (.Y(N5554), .A0(N18501), .A1(N18439), .B0(N18249), .B1(N18933));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4134 (.Y(N5555), .A(N18510), .B(N18573));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4135 (.Y(N5558), .A0(N18510), .A1(N18398), .B0(N18420), .B1(N18933));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4138 (.Y(N18335), .A0(N18510), .A1(N18572), .B0(N18901), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4139 (.Y(N18337), .A0(N18510), .A1(N18430), .B0(N18889), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4141 (.Y(N18339), .A0(N18510), .A1(N18901), .B0(N18448), .B1(N18933));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I4142 (.Y(N18341), .A(N18510), .B(N18405));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4150 (.Y(N5578), .A(N18510), .B(N18476));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4152 (.Y(N5584), .A0(N18510), .A1(N18249), .B0(N18405), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4153 (.Y(N18343), .A0(N18510), .A1(N18901), .B0(N18439), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4154 (.Y(N5586), .A0(N18510), .A1(N18572), .B0(N18448), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4157 (.Y(N5591), .A0(N18510), .A1(N18249), .B0(N18439), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4158 (.Y(N5592), .A0(N18510), .A1(N18889), .B0(N18901), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4159 (.Y(N5593), .A0(N18510), .A1(N18249), .B0(N18470), .B1(N18933));
INVXL inst_noninc_a_cellmath__55_2WWMM_I4160 (.Y(N5594), .A(N18460));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I14513 (.Y(N18820), .A0(N18933), .A1(N18572), .B0(N18889), .B1(N18510));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4164 (.Y(N18347), .A0(N18510), .A1(N18409), .B0(N18460), .B1(N18933));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I4933 (.Y(N6610), .A0(N18510), .A1(N18410), .B0(N18477), .B1(N18933));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I4934 (.Y(N18349), .A0(N18510), .A1(N18410), .B0(N18405), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4936 (.Y(N6613), .A0(N18510), .A1(N18399), .B0(N18458), .B1(N18933));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I4949 (.Y(N6633), .A(N18510), .B(N18572));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I4950 (.Y(N6635), .A(N18249), .B(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4952 (.Y(N6638), .A0(N18510), .A1(N18470), .B0(N18409), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4955 (.Y(N6641), .A0(N18514), .A1(N18470), .B0(N18249), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4956 (.Y(N6642), .A0(N18514), .A1(N18572), .B0(N18409), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4957 (.Y(N6643), .A0(N18514), .A1(N18405), .B0(N18458), .B1(N18937));
INVXL inst_noninc_a_cellmath__55_2WWMM_I4961 (.Y(N6648), .A(N18448));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4963 (.Y(N18351), .A(N18514), .B(N18897));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4965 (.Y(N18353), .A0(N18399), .A1(N18514), .B0(N18410), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4966 (.Y(N6657), .A0(N18510), .A1(N18405), .B0(N18249), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I14516 (.Y(N18831), .A0(N18937), .A1(N18430), .B0(N18510), .B1(N18889));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4975 (.Y(N6670), .A0(N18677), .A1(N18337), .B0(N18331), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4976 (.Y(N6671), .A0(N18677), .A1(N4351), .B0(N18259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4977 (.Y(N6672), .A0(N18677), .A1(N18311), .B0(N5537), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4978 (.Y(N6673), .A0(N18677), .A1(N18343), .B0(N18735), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4985 (.Y(N6683), .A0(N18677), .A1(N18281), .B0(N5550), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4986 (.Y(N6684), .A0(N18677), .A1(N1103), .B0(N18748), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4987 (.Y(N6685), .A0(N18677), .A1(N6610), .B0(N18333), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I4988 (.Y(N6686), .A0(N18677), .A1(N18349), .B0(N5553), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4989 (.Y(N6687), .A(N18672), .B(N5554));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4990 (.Y(N6690), .A0(N18672), .A1(N6613), .B0(N5555), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4991 (.Y(N6691), .A0(N18672), .A1(N18546), .B0(N5558), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4992 (.Y(N6692), .A0(N18672), .A1(N18889), .B0(N18735), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4993 (.Y(N6693), .A0(N18672), .A1(N18407), .B0(N18277), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4994 (.Y(N6694), .A0(N18677), .A1(N18265), .B0(N18335), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4995 (.Y(N6695), .A0(N18677), .A1(N18311), .B0(N18337), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4996 (.Y(N6696), .A0(N18677), .A1(N18335), .B0(N18275), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4997 (.Y(N6697), .A0(N18677), .A1(N18315), .B0(N18339), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4998 (.Y(N6698), .A0(N18677), .A1(N18596), .B0(N18341), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5003 (.Y(N6707), .A0(N18677), .A1(N6633), .B0(N18739), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5004 (.Y(N6708), .A0(N18677), .A1(N6635), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5005 (.Y(N6709), .A0(N18677), .A1(N18287), .B0(N18265), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5006 (.Y(N6710), .A0(N18677), .A1(N6638), .B0(N5578), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5007 (.Y(N6711), .A0(N18677), .A1(N18297), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5008 (.Y(N6712), .A0(N18672), .A1(N18333), .B0(N5584), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5009 (.Y(N6713), .A0(N18672), .A1(N6641), .B0(N18343), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5010 (.Y(N6714), .A0(N18672), .A1(N6642), .B0(N5586), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5011 (.Y(N6715), .A0(N18672), .A1(N6643), .B0(N2163), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5012 (.Y(N6716), .A0(N18672), .A1(N5591), .B0(N18341), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5013 (.Y(N6717), .A0(N18672), .A1(N18235), .B0(N5591), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5014 (.Y(N6718), .A0(N18672), .A1(N18341), .B0(N5592), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5015 (.Y(N6719), .A0(N18672), .A1(N6648), .B0(N5593), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5016 (.Y(N6720), .A0(N18672), .A1(N2163), .B0(N5594), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5017 (.Y(N6721), .A0(N18672), .A1(N18351), .B0(N18820), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5018 (.Y(N6722), .A0(N18672), .A1(N18583), .B0(N18609), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5019 (.Y(N6723), .A0(N18672), .A1(N18353), .B0(N18730), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5020 (.Y(N6724), .A0(N6657), .A1(N18672), .B0(N18347), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5021 (.Y(N6725), .A0(N18672), .A1(N18831), .B0(N18729), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5022 (.Y(N6726), .A0(N18672), .A1(N18735), .B0(N18601), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5023 (.Y(N6727), .A0(N18247), .A1(N18677), .B0(N18323), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I5778 (.Y(N7736), .A(N18439), .B(N18937));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I5779 (.Y(N18357), .A0(N18510), .A1(N18399), .B0(N18430), .B1(N18933));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14161 (.Y(N18832), .A(N18357));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14163 (.Y(N18834), .A(N18832));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14162 (.Y(N18833), .A(N18832));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5780 (.Y(N7739), .A0(N18510), .A1(N18573), .B0(N18420), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5787 (.Y(N7753), .A0(N18510), .A1(N18439), .B0(N18889), .B1(N18933));
INVXL inst_noninc_a_cellmath__55_2WWMM_I5789 (.Y(N7755), .A(N18249));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5793 (.Y(N7759), .A0(N18514), .A1(N18470), .B0(N18572), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5806 (.Y(N7780), .A0(N18514), .A1(N18889), .B0(N18477), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5808 (.Y(N7783), .A0(N18514), .A1(N18430), .B0(N18458), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5815 (.Y(N7790), .A0(N18514), .A1(N18405), .B0(N18448), .B1(N18933));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I5820 (.Y(N7795), .A(N18514), .B(N18418));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5823 (.Y(N7799), .A0(N18514), .A1(N18477), .B0(N18399), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6579 (.Y(N8814), .A0(N18514), .A1(N18477), .B0(N18418), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6581 (.Y(N18359), .A0(N18514), .A1(N18573), .B0(N18399), .B1(N18933));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I6583 (.Y(N8819), .A0(N18514), .A1(N18448), .B0(N18439), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6590 (.Y(N8831), .A0(N18514), .A1(N18470), .B0(N18458), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6597 (.Y(N8843), .A0(N18514), .A1(N18458), .B0(N18897), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6599 (.Y(N8845), .A0(N18514), .A1(N18410), .B0(N18889), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6608 (.Y(N8861), .A0(N18514), .A1(N18430), .B0(N18897), .B1(N18933));
INVXL inst_noninc_a_cellmath__55_2WWMM_I6609 (.Y(N8862), .A(N18478));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6610 (.Y(N8863), .A(N18430), .B(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6613 (.Y(N8867), .A0(N18514), .A1(N18470), .B0(N18439), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6614 (.Y(N8868), .A0(N18514), .A1(N18458), .B0(N18470), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6616 (.Y(N8870), .A0(N18514), .A1(N18430), .B0(N18410), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6617 (.Y(N8871), .A0(N18514), .A1(N18439), .B0(N18410), .B1(N18933));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6619 (.Y(N8873), .A(N18937), .B(N18399));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6624 (.Y(N18361), .A0(N18514), .A1(N18450), .B0(N18897), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6633 (.Y(N8895), .A0(N18677), .A1(N8814), .B0(N18327), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6634 (.Y(N8896), .A0(N18677), .A1(N18341), .B0(N7736), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6635 (.Y(N8897), .A0(N18677), .A1(N18359), .B0(N18834), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6636 (.Y(N8898), .A0(N18677), .A1(N18319), .B0(N7739), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6637 (.Y(N8899), .A0(N18677), .A1(N8819), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6638 (.Y(N8900), .A0(N18677), .A1(N18231), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6639 (.Y(N8901), .A(N18301), .B(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6643 (.Y(N8909), .A0(N18677), .A1(N6610), .B0(N7753), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6644 (.Y(N8910), .A0(N18677), .A1(N8831), .B0(N18337), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6645 (.Y(N8911), .A0(N18672), .A1(N5578), .B0(N7755), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6646 (.Y(N8912), .A0(N18672), .A1(N5558), .B0(N2180), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6647 (.Y(N8913), .A0(N18672), .A1(N5578), .B0(N18748), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6648 (.Y(N8914), .A0(N18672), .A1(N4371), .B0(N2179), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6649 (.Y(N8915), .A0(N18672), .A1(N2175), .B0(N7759), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6650 (.Y(N8916), .A0(N18672), .A1(N18609), .B0(N7736), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6651 (.Y(N8917), .A(N18672), .B(N8843));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6652 (.Y(N8919), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18579));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6653 (.Y(N8922), .A0(N18672), .A1(N8845), .B0(N18399), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6654 (.Y(N8923), .A0(N18672), .A1(N18319), .B0(N18569), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6655 (.Y(N8924), .A0(N18672), .A1(N18601), .B0(N18265), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6656 (.Y(N8925), .A0(N18672), .A1(N18247), .B0(N18269), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6657 (.Y(N8926), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B(N18341));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6661 (.Y(N8933), .A0(N18672), .A1(N18327), .B0(N1068), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6662 (.Y(N8934), .A0(N18672), .A1(N8861), .B0(N7780), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6663 (.Y(N8935), .A0(N18672), .A1(N8862), .B0(N18514), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6664 (.Y(N8936), .A0(N18672), .A1(N8863), .B0(N7783), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6665 (.Y(N8937), .A0(N18677), .A1(N1086), .B0(N18321), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6666 (.Y(N8938), .A0(N18677), .A1(N18706), .B0(N6638), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6667 (.Y(N8939), .A0(N18677), .A1(N8867), .B0(N5592), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6668 (.Y(N8940), .A0(N18677), .A1(N8868), .B0(N18331), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6669 (.Y(N8941), .A0(N18677), .A1(N18353), .B0(N18275), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6670 (.Y(N8942), .A0(N18677), .A1(N8870), .B0(N18277), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6671 (.Y(N8943), .A0(N18677), .A1(N8871), .B0(N7790), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6672 (.Y(N8944), .A0(N18677), .A1(N18337), .B0(N18579), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6673 (.Y(N8945), .A0(N18677), .A1(N8873), .B0(N1066), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6674 (.Y(N8946), .A0(N18677), .A1(N18331), .B0(N18273), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6675 (.Y(N8947), .A0(N18672), .A1(N6635), .B0(N18297), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6676 (.Y(N8948), .A0(N18672), .A1(N18831), .B0(N7795), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6677 (.Y(N8949), .A0(N18672), .A1(N18347), .B0(N18291), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6678 (.Y(N8950), .A0(N18672), .A1(N18361), .B0(N18349), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6679 (.Y(N8951), .A0(N18672), .A1(N18353), .B0(N7799), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6680 (.Y(N8952), .A0(N18672), .A1(N7739), .B0(N18275), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6681 (.Y(N8953), .A0(N18672), .A1(N18301), .B0(N18253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6682 (.Y(N8954), .A0(N18672), .A1(N18231), .B0(N18253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6687 (.Y(N8962), .A0(N18802), .A1(N8895), .B0(N6670), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6688 (.Y(N8963), .A0(N18802), .A1(N8896), .B0(N6671), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6689 (.Y(N8964), .A0(N18802), .A1(N8897), .B0(N6672), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6690 (.Y(N8965), .A0(N18802), .A1(N8898), .B0(N6673), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6691 (.Y(N8966), .A0(N18802), .A1(N8899), .B0(N4469), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6692 (.Y(N8967), .A0(N18802), .A1(N8900), .B0(N4473), .B1(N19085));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6693 (.Y(N8968), .A(N18802), .B(N8901));
NOR2XL andori2bb1_A_I14587 (.Y(N19132), .A(N18677), .B(N18231));
NOR2XL andori2bb1_A_I14588 (.Y(N8972), .A(N19132), .B(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6697 (.Y(N8977), .A0(N18802), .A1(N8909), .B0(N6683), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6698 (.Y(N8978), .A0(N18802), .A1(N8910), .B0(N6684), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6699 (.Y(N8979), .A0(N18802), .A1(N8911), .B0(N6685), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6700 (.Y(N8980), .A0(N18802), .A1(N8912), .B0(N6686), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6701 (.Y(N8981), .A0(N18802), .A1(N8913), .B0(N6687), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6702 (.Y(N8982), .A0(N18802), .A1(N8914), .B0(N6690), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6703 (.Y(N8983), .A0(N18802), .A1(N8915), .B0(N6691), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6704 (.Y(N8984), .A0(N18802), .A1(N8916), .B0(N6692), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6705 (.Y(N8985), .A0(N18802), .A1(N8917), .B0(N6693), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6706 (.Y(N8986), .A0(N18802), .A1(N8919), .B0(N6694), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6707 (.Y(N8987), .A0(N18802), .A1(N8922), .B0(N6695), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6708 (.Y(N8988), .A0(N18802), .A1(N8923), .B0(N6696), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6709 (.Y(N8989), .A0(N18802), .A1(N8924), .B0(N6697), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6710 (.Y(N8990), .A0(N18802), .A1(N8925), .B0(N6698), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6711 (.Y(N8991), .A0(N18802), .A1(N8926), .B0(N2261), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6715 (.Y(N8998), .A0(N18802), .A1(N8933), .B0(N6707), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6716 (.Y(N8999), .A0(N18802), .A1(N8934), .B0(N6708), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6717 (.Y(N9000), .A0(N18802), .A1(N8935), .B0(N6709), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6718 (.Y(N9001), .A0(N18802), .A1(N8936), .B0(N6710), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6719 (.Y(N9002), .A0(N18802), .A1(N8937), .B0(N6711), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6720 (.Y(N9003), .A0(N18802), .A1(N8938), .B0(N6712), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6721 (.Y(N9004), .A0(N18802), .A1(N8939), .B0(N6713), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6722 (.Y(N9005), .A0(N18802), .A1(N8940), .B0(N6714), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6723 (.Y(N9006), .A0(N18802), .A1(N8941), .B0(N6715), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6724 (.Y(N9007), .A0(N18802), .A1(N8942), .B0(N6716), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6725 (.Y(N9008), .A0(N18802), .A1(N8943), .B0(N6717), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6726 (.Y(N9009), .A0(N18802), .A1(N8944), .B0(N6718), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6727 (.Y(N9010), .A0(N18802), .A1(N8945), .B0(N6719), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6728 (.Y(N9011), .A0(N18802), .A1(N8946), .B0(N6720), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6729 (.Y(N9012), .A0(N18802), .A1(N8947), .B0(N6721), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6730 (.Y(N9013), .A0(N18802), .A1(N8948), .B0(N6722), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6731 (.Y(N9014), .A0(N18802), .A1(N8949), .B0(N6723), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6732 (.Y(N9015), .A0(N18802), .A1(N8950), .B0(N6724), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6733 (.Y(N9016), .A0(N18802), .A1(N8951), .B0(N6725), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6734 (.Y(N9017), .A0(N18802), .A1(N8952), .B0(N6726), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6735 (.Y(N9018), .A0(N18802), .A1(N8953), .B0(N6727), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6736 (.Y(N9019), .A0(N18802), .A1(N8954), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B1(N19086));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I14519 (.Y(N9020), .A0N(N18253), .A1N(inst_noninc_a_cellmath__55_2WWMM_in0[19]), .B0(N18802));
NOR2XL andori2bb1_A_I14589 (.Y(N19139), .A(N18672), .B(N18323));
NOR2XL andori2bb1_A_I14590 (.Y(N9022), .A(N19139), .B(N19086));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14531 (.Y(N19107), .A(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14441 (.Y(N19112), .A(N19107));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14194 (.Y(N18865), .A(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6741 (.Y(N9028), .A0(N18865), .A1(N8962), .B0(N4478), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6742 (.Y(N9029), .A0(N18865), .A1(N8963), .B0(N4479), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6743 (.Y(N9030), .A0(N18865), .A1(N8964), .B0(N4480), .B1(N19112));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14440 (.Y(N19111), .A(N19107));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6744 (.Y(N9031), .A0(N18865), .A1(N8965), .B0(N4481), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6745 (.Y(N9032), .A0(N18865), .A1(N8966), .B0(N4482), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6746 (.Y(N9033), .A0(N18865), .A1(N8967), .B0(N4483), .B1(N19111));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6747 (.Y(N9034), .A(N18865), .B(N8968));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6748 (.Y(N9036), .A(N19111), .B(N8968));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6749 (.Y(N9039), .A(N18865), .B(N8972));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6751 (.Y(N9042), .A0(N18865), .A1(N8977), .B0(N4493), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6752 (.Y(N9043), .A0(N18865), .A1(N8978), .B0(N4494), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6753 (.Y(N9044), .A0(N18865), .A1(N8979), .B0(N4495), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6754 (.Y(N9045), .A0(N18865), .A1(N8980), .B0(N4496), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6755 (.Y(N9046), .A0(N18865), .A1(N8981), .B0(N4497), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6756 (.Y(N9047), .A0(N18865), .A1(N8982), .B0(N4498), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6757 (.Y(N9048), .A0(N18865), .A1(N8983), .B0(N4499), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6758 (.Y(N9049), .A0(N18865), .A1(N8984), .B0(N4500), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6759 (.Y(N9050), .A0(N18865), .A1(N8985), .B0(N4501), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6760 (.Y(N9051), .A0(N18865), .A1(N8986), .B0(N4502), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6761 (.Y(N9052), .A0(N18865), .A1(N8987), .B0(N4503), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6762 (.Y(N9053), .A0(N18865), .A1(N8988), .B0(N4504), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6763 (.Y(N9054), .A0(N18865), .A1(N8989), .B0(N4505), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6764 (.Y(N9055), .A0(N18865), .A1(N8990), .B0(N4506), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6765 (.Y(N9056), .A0(N18865), .A1(N8991), .B0(N4507), .B1(N19111));
NOR2XL andori2bb1_A_I14591 (.Y(N19146), .A(N18802), .B(N18283));
NOR2XL andori2bb1_A_I14592 (.Y(N9057), .A(N19146), .B(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6769 (.Y(N9063), .A0(N18865), .A1(N8998), .B0(N4513), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6770 (.Y(N9064), .A0(N18865), .A1(N8999), .B0(N4514), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6771 (.Y(N9065), .A0(N18865), .A1(N9000), .B0(N4515), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6772 (.Y(N9066), .A0(N18865), .A1(N9001), .B0(N4516), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6773 (.Y(N9067), .A0(N18865), .A1(N9002), .B0(N4517), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6774 (.Y(N9068), .A0(N18865), .A1(N9003), .B0(N4518), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6775 (.Y(N9069), .A0(N18865), .A1(N9004), .B0(N4519), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6776 (.Y(N9070), .A0(N18865), .A1(N9005), .B0(N4520), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6777 (.Y(N9071), .A0(N18865), .A1(N9006), .B0(N4521), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6778 (.Y(N9072), .A0(N18865), .A1(N9007), .B0(N4522), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6779 (.Y(N9073), .A0(N18865), .A1(N9008), .B0(N4523), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6780 (.Y(N9074), .A0(N18865), .A1(N9009), .B0(N4524), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6781 (.Y(N9075), .A0(N18865), .A1(N9010), .B0(N4525), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6782 (.Y(N9076), .A0(N18865), .A1(N9011), .B0(N4526), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6783 (.Y(N9077), .A0(N18865), .A1(N9012), .B0(N4527), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6784 (.Y(N9078), .A0(N18865), .A1(N9013), .B0(N4528), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6785 (.Y(N9079), .A0(N18865), .A1(N9014), .B0(N4529), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6786 (.Y(N9080), .A0(N18865), .A1(N9015), .B0(N4530), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6787 (.Y(N9081), .A0(N18865), .A1(N9016), .B0(N4531), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6788 (.Y(N9082), .A0(N18865), .A1(N9017), .B0(N4532), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6789 (.Y(N9083), .A0(N18865), .A1(N9018), .B0(N4533), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6790 (.Y(N9084), .A0(N18865), .A1(N9019), .B0(N4534), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6791 (.Y(N9085), .A0(N18865), .A1(N9020), .B0(N4535), .B1(N19112));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6792 (.Y(N9086), .A(N18865), .B(N9022));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7559 (.Y(N10112), .A0(N18514), .A1(N18399), .B0(N18897), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7575 (.Y(N10134), .A0(N18531), .A1(N18573), .B0(N18458), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7577 (.Y(N10137), .A0(N18531), .A1(N18458), .B0(N18405), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7584 (.Y(N10146), .A0(N18531), .A1(N18418), .B0(N18399), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8348 (.Y(N11159), .A0(N18531), .A1(N18249), .B0(N18573), .B1(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8361 (.Y(N11176), .A(N18405), .B(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I8362 (.Y(N11178), .A(N18531), .B(N18400));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8363 (.Y(N11181), .A(N18573), .B(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8377 (.Y(N11204), .A0(N18531), .A1(N18418), .B0(N18450), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8379 (.Y(N11207), .A0(N18531), .A1(N18450), .B0(N18470), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8382 (.Y(N11210), .A0(N18531), .A1(N18897), .B0(N18249), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8399 (.Y(N11236), .A0(N18672), .A1(N18341), .B0(N7799), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8400 (.Y(N11237), .A0(N18677), .A1(N18359), .B0(N3314), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8401 (.Y(N11238), .A0(N18677), .A1(N18229), .B0(N18259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8402 (.Y(N11239), .A0(N18677), .A1(N11159), .B0(N5537), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8403 (.Y(N11240), .A0(N18677), .A1(N7790), .B0(N18601), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8404 (.Y(N11241), .A0(N18677), .A1(N18546), .B0(N18253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8405 (.Y(N11242), .A0(N18672), .A1(N18341), .B0(N18323), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8406 (.Y(N11243), .A(N18672), .B(N18247));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8409 (.Y(N11248), .A0(N18672), .A1(N1084), .B0(N18343), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8410 (.Y(N11249), .A0(N18672), .A1(N6641), .B0(N4342), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8411 (.Y(N11250), .A0(N18672), .A1(N18233), .B0(N18297), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8412 (.Y(N11251), .A0(N18672), .A1(N5558), .B0(N18833), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8413 (.Y(N11252), .A0(N18672), .A1(N4377), .B0(N4367), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8414 (.Y(N11253), .A0(N18672), .A1(N4377), .B0(N5554), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8415 (.Y(N11254), .A0(N18672), .A1(N11176), .B0(N10112), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8416 (.Y(N11255), .A0(N18672), .A1(N11178), .B0(N18341), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8417 (.Y(N11256), .A0(N18672), .A1(N11181), .B0(N18399), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8418 (.Y(N11257), .A0(N18672), .A1(N18833), .B0(N18569), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8419 (.Y(N11258), .A0(N18672), .A1(N18569), .B0(N18748), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8420 (.Y(N11259), .A0(N18672), .A1(N18321), .B0(N18609), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8427 (.Y(N11271), .A0(N18672), .A1(N8861), .B0(N18339), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8428 (.Y(N11272), .A0(N18672), .A1(N3314), .B0(N18291), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8429 (.Y(N11273), .A0(N18672), .A1(N18353), .B0(N18307), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8430 (.Y(N11274), .A0(N18672), .A1(N18247), .B0(N10112), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8431 (.Y(N11275), .A0(N18672), .A1(N11204), .B0(N10134), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8432 (.Y(N11276), .A0(N18672), .A1(N18908), .B0(N18889), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8433 (.Y(N11277), .A0(N18672), .A1(N11207), .B0(N10137), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8434 (.Y(N11278), .A0(N18672), .A1(N11207), .B0(N8862), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8435 (.Y(N11279), .A0(N18672), .A1(N18321), .B0(N3306), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8436 (.Y(N11280), .A0(N18672), .A1(N11210), .B0(N18273), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8437 (.Y(N11281), .A0(N18672), .A1(N18531), .B0(N18243), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8438 (.Y(N11282), .A0(N18677), .A1(N5550), .B0(N18729), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8439 (.Y(N11283), .A0(N18677), .A1(N18259), .B0(N18725), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8440 (.Y(N11284), .A0(N18677), .A1(N5553), .B0(N10146), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8441 (.Y(N11285), .A0(N18677), .A1(N2140), .B0(N18820), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8442 (.Y(N11286), .A0(N18677), .A1(N18596), .B0(N18609), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8443 (.Y(N11287), .A(N18361), .B(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8445 (.Y(N11292), .A0(N18677), .A1(N18400), .B0(N18820), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8446 (.Y(N11293), .A0(N18677), .A1(N18897), .B0(N7790), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8447 (.Y(N11294), .A0(N18677), .A1(N1102), .B0(N18546), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8448 (.Y(N11295), .A0(N18677), .A1(N18247), .B0(N18341), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I8449 (.Y(N11296), .A(N18677), .B(N18247));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I9211 (.Y(N12316), .A(N18889), .B(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I9213 (.Y(N12319), .A0(N18531), .A1(N18478), .B0(N18889), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9218 (.Y(N12328), .A0(N18531), .A1(N18405), .B0(N18430), .B1(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I9229 (.Y(N12343), .A(N18531), .B(N18430));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9230 (.Y(N12346), .A0(N18531), .A1(N18450), .B0(N18889), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9237 (.Y(N12357), .A0(N18531), .A1(N18430), .B0(N18470), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9240 (.Y(N12362), .A0(N18531), .A1(N18430), .B0(N18450), .B1(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I9241 (.Y(N12363), .A(N18531), .B(N18458));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9242 (.Y(N12366), .A0(N18531), .A1(N18418), .B0(N18411), .B1(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I9243 (.Y(N12367), .A(N18458), .B(N18937));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10013 (.Y(N13404), .A(N18531), .B(N18460));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10014 (.Y(N13406), .A0(N18531), .A1(N18885), .B0(N18405), .B1(N18937));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I10015 (.Y(N13407), .A0(N18531), .A1(N18478), .B0(N18249), .B1(N18937));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I10016 (.Y(N13408), .A(N18531), .B(N18411));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10017 (.Y(N13411), .A0(N18531), .A1(N18420), .B0(N18430), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10032 (.Y(N13437), .A0(N18531), .A1(N18405), .B0(N18478), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10036 (.Y(N13443), .A0(N18531), .A1(N18460), .B0(N18450), .B1(N18937));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10040 (.Y(N13448), .A0(N18531), .A1(N18430), .B0(N18420), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10048 (.Y(N13459), .A0(N18531), .A1(N18411), .B0(N18470), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10051 (.Y(N13462), .A0(N18531), .A1(N18420), .B0(N18439), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10057 (.Y(N13471), .A0(N18677), .A1(N1044), .B0(N4350), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10058 (.Y(N13472), .A0(N18677), .A1(N7739), .B0(N18351), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10059 (.Y(N13473), .A0(N18677), .A1(N18231), .B0(N18702), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I10062 (.Y(N13477), .A(N18281));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10063 (.Y(N13478), .A0(N18677), .A1(N18269), .B0(N18596), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10067 (.Y(N13487), .A0(N18677), .A1(N13404), .B0(N12316), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10068 (.Y(N13488), .A0(N18677), .A1(N13406), .B0(N18717), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I10069 (.Y(N13489), .A0(N18677), .A1(N13407), .B0(N12319), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10070 (.Y(N13490), .A0(N13408), .A1(N18677), .B0(N18347), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10071 (.Y(N13491), .A0(N18677), .A1(N13411), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10072 (.Y(N13492), .A0(N18677), .A1(N18331), .B0(N18351), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10073 (.Y(N13493), .A0(N18677), .A1(N18353), .B0(N4380), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10074 (.Y(N13494), .A0(N18677), .A1(N5554), .B0(N12328), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10075 (.Y(N13495), .A0(N18677), .A1(N12343), .B0(N18293), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10076 (.Y(N13496), .A0(N18677), .A1(N18253), .B0(N18295), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10077 (.Y(N13497), .A0(N18677), .A1(N18323), .B0(N4351), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10078 (.Y(N13498), .A0(N18677), .A1(N18885), .B0(N6610), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10079 (.Y(N13499), .A0(N18677), .A1(N18405), .B0(N2180), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10081 (.Y(N13501), .A0(N18677), .A1(N18247), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10085 (.Y(N13508), .A0(N18677), .A1(N2142), .B0(N12343), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10086 (.Y(N13509), .A0(N18677), .A1(N13437), .B0(N12346), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10087 (.Y(N13510), .A0(N18677), .A1(N2147), .B0(N12343), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10088 (.Y(N13511), .A0(N18677), .A1(N18333), .B0(N18359), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10089 (.Y(N13512), .A0(N18677), .A1(N18253), .B0(N18820), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10090 (.Y(N13513), .A0(N18677), .A1(N13443), .B0(N18735), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10091 (.Y(N13514), .A0(N18677), .A1(N12367), .B0(N7783), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10092 (.Y(N13515), .A0(N18672), .A1(N7799), .B0(N3309), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10093 (.Y(N13516), .A0(N18672), .A1(N1084), .B0(N12357), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10094 (.Y(N13517), .A0(N18672), .A1(N13448), .B0(N3306), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10095 (.Y(N13518), .A0(N18672), .A1(N18339), .B0(N18361), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10096 (.Y(N13519), .A0(N18672), .A1(N18546), .B0(N12362), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10097 (.Y(N13520), .A0(N18672), .A1(N18407), .B0(N12363), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10098 (.Y(N13521), .A0(N18672), .A1(N6642), .B0(N12366), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10099 (.Y(N13522), .A0(N18672), .A1(N18351), .B0(N12367), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10100 (.Y(N13523), .A0(N18672), .A1(N12367), .B0(N18820), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10101 (.Y(N13524), .A0(N18672), .A1(N18353), .B0(N18343), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10102 (.Y(N13525), .A0(N18677), .A1(N13459), .B0(N18908), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10103 (.Y(N13526), .A0(N18677), .A1(N18748), .B0(N4329), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10104 (.Y(N13527), .A0(N18677), .A1(N18725), .B0(N18293), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10105 (.Y(N13528), .A0(N18677), .A1(N13462), .B0(N18361), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10106 (.Y(N13529), .A0(N18677), .A1(N18531), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10111 (.Y(N13538), .A0(N18802), .A1(N13471), .B0(N11236), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10112 (.Y(N13539), .A0(N18802), .A1(N13472), .B0(N11237), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10113 (.Y(N13540), .A0(N18802), .A1(N13473), .B0(N11238), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10114 (.Y(N13541), .A0(N18802), .A1(N18400), .B0(N11239), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10115 (.Y(N13542), .A0(N18802), .A1(N18411), .B0(N11240), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10116 (.Y(N13543), .A0(N18802), .A1(N13477), .B0(N11241), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10117 (.Y(N13544), .A0(N18802), .A1(N13478), .B0(N11242), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10118 (.Y(N13545), .A0(N18802), .A1(N18283), .B0(N11243), .B1(N19085));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10119 (.Y(N13546), .A(N18802), .B(N18283));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10121 (.Y(N13551), .A0(N18802), .A1(N13487), .B0(N11248), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10122 (.Y(N13552), .A0(N18802), .A1(N13488), .B0(N11249), .B1(N19085));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I10123 (.Y(N13553), .A0(N18802), .A1(N13489), .B0(N11250), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10124 (.Y(N13554), .A0(N18802), .A1(N13490), .B0(N11251), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10125 (.Y(N13555), .A0(N18802), .A1(N13491), .B0(N11252), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10126 (.Y(N13556), .A0(N18802), .A1(N13492), .B0(N11253), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10127 (.Y(N13557), .A0(N18802), .A1(N13493), .B0(N11254), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10128 (.Y(N13558), .A0(N18802), .A1(N13494), .B0(N11255), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10129 (.Y(N13559), .A0(N18802), .A1(N13495), .B0(N11256), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10130 (.Y(N13560), .A0(N18802), .A1(N13496), .B0(N11257), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10131 (.Y(N13561), .A0(N18802), .A1(N13497), .B0(N11258), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10132 (.Y(N13562), .A0(N18802), .A1(N13498), .B0(N11259), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10133 (.Y(N13563), .A0(N18802), .A1(N13499), .B0(N4436), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10134 (.Y(N13564), .A0(N18802), .A1(N2202), .B0(N4437), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10135 (.Y(N13565), .A0(N18802), .A1(N13501), .B0(N18329), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10136 (.Y(N13566), .A0(N18802), .A1(N8926), .B0(N18329), .B1(N19085));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10137 (.Y(N13567), .A(N18329), .B(N19085));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I10138 (.Y(N13569), .A(N18802), .B(N2253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10139 (.Y(N13572), .A0(N18802), .A1(N13508), .B0(N11271), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10140 (.Y(N13573), .A0(N18802), .A1(N13509), .B0(N11272), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10141 (.Y(N13574), .A0(N18802), .A1(N13510), .B0(N11273), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10142 (.Y(N13575), .A0(N18802), .A1(N13511), .B0(N11274), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10143 (.Y(N13576), .A0(N18802), .A1(N13512), .B0(N11275), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10144 (.Y(N13577), .A0(N18802), .A1(N13513), .B0(N11276), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10145 (.Y(N13578), .A0(N18802), .A1(N13514), .B0(N11277), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10146 (.Y(N13579), .A0(N18802), .A1(N13515), .B0(N11278), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10147 (.Y(N13580), .A0(N18802), .A1(N13516), .B0(N11279), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10148 (.Y(N13581), .A0(N18802), .A1(N13517), .B0(N11280), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10149 (.Y(N13582), .A0(N18802), .A1(N13518), .B0(N11281), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10150 (.Y(N13583), .A0(N18802), .A1(N13519), .B0(N11282), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10151 (.Y(N13584), .A0(N18802), .A1(N13520), .B0(N11283), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10152 (.Y(N13585), .A0(N18802), .A1(N13521), .B0(N11284), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10153 (.Y(N13586), .A0(N18802), .A1(N13522), .B0(N11285), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10154 (.Y(N13587), .A0(N18802), .A1(N13523), .B0(N11286), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10155 (.Y(N13588), .A0(N18802), .A1(N13524), .B0(N11287), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10156 (.Y(N13589), .A0(N18802), .A1(N13525), .B0(N4417), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10157 (.Y(N13590), .A0(N18802), .A1(N13526), .B0(N11292), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10158 (.Y(N13591), .A0(N18802), .A1(N13527), .B0(N11293), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10159 (.Y(N13592), .A0(N18802), .A1(N13528), .B0(N11294), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10160 (.Y(N13593), .A0(N18802), .A1(N13529), .B0(N11295), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10161 (.Y(N13594), .A0(N18802), .A1(N8901), .B0(N11296), .B1(N19085));
INVXL inst_noninc_a_cellmath__55_2WWMM_I10923 (.Y(N14617), .A(N18440));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I10925 (.Y(N14619), .A0(N18531), .A1(N18440), .B0(N18478), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10927 (.Y(N14621), .A0(N18531), .A1(N18897), .B0(N18420), .B1(N18933));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10941 (.Y(N14638), .A0(N18531), .A1(N18897), .B0(N18400), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10944 (.Y(N14641), .A0(N18531), .A1(N18885), .B0(N18450), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10950 (.Y(N14649), .A0(N18531), .A1(N18430), .B0(N18249), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10956 (.Y(N14658), .A0(N18531), .A1(N18400), .B0(N18478), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11728 (.Y(N15695), .A0(N18531), .A1(N18479), .B0(N18470), .B1(N18909));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14240 (.Y(N18911), .A(N18907));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11738 (.Y(N15708), .A0(N18531), .A1(N18470), .B0(N18450), .B1(N18911));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11750 (.Y(N15724), .A0(N18531), .A1(N18460), .B0(N18420), .B1(N18911));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11751 (.Y(N15725), .A0(N18531), .A1(N18450), .B0(N18479), .B1(N18911));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11769 (.Y(N15750), .A0(N18677), .A1(N18706), .B0(N8868), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11770 (.Y(N15751), .A0(N18677), .A1(N5592), .B0(N6657), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11771 (.Y(N15752), .A0(N18677), .A1(N18722), .B0(N18831), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11772 (.Y(N15753), .A0(N18677), .A1(N7759), .B0(N18259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11773 (.Y(N15754), .A0(N18677), .A1(N18277), .B0(N18706), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11774 (.Y(N15755), .A0(N18677), .A1(N18349), .B0(N18361), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11775 (.Y(N15756), .A0(N18677), .A1(N18315), .B0(N18231), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11779 (.Y(N15762), .A0(N18677), .A1(N4342), .B0(N14617), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11780 (.Y(N15763), .A0(N18677), .A1(N18259), .B0(N18287), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11781 (.Y(N15764), .A0(N18677), .A1(N4344), .B0(N14619), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11782 (.Y(N15765), .A0(N18672), .A1(N15695), .B0(N8819), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11783 (.Y(N15766), .A0(N18672), .A1(N18335), .B0(N14621), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11784 (.Y(N15767), .A0(N18672), .A1(N4344), .B0(N8867), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11785 (.Y(N15768), .A0(N18672), .A1(N18729), .B0(N13448), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11786 (.Y(N15769), .A0(N18672), .A1(N8873), .B0(N2175), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I11787 (.Y(N15770), .A0(N4371), .A1(N18677), .B0(N18609), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11788 (.Y(N15771), .A0(N18677), .A1(N8845), .B0(N8843), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11789 (.Y(N15772), .A0(N18677), .A1(N18319), .B0(N18579), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11790 (.Y(N15773), .A0(N18677), .A1(N18259), .B0(N18359), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11791 (.Y(N15774), .A0(N18677), .A1(N18729), .B0(N8861), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11792 (.Y(N15775), .A0(N18677), .A1(N15708), .B0(N18579), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11793 (.Y(N15776), .A0(N18677), .A1(N18531), .B0(N18341), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11797 (.Y(N15783), .A0(N18677), .A1(N8845), .B0(N14638), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11798 (.Y(N15784), .A0(N18677), .A1(N18339), .B0(N18261), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11799 (.Y(N15785), .A0(N18677), .A1(N8831), .B0(N18339), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11800 (.Y(N15786), .A0(N18672), .A1(N18729), .B0(N14641), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11801 (.Y(N15787), .A0(N18672), .A1(N18831), .B0(N5555), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11802 (.Y(N15788), .A0(N18672), .A1(N15708), .B0(N18277), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11803 (.Y(N15789), .A0(N18672), .A1(N18748), .B0(N18333), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11804 (.Y(N15790), .A0(N18672), .A1(N15724), .B0(N18349), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11805 (.Y(N15791), .A0(N18672), .A1(N15725), .B0(N18235), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11806 (.Y(N15792), .A0(N18672), .A1(N15724), .B0(N14649), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11807 (.Y(N15793), .A0(N18672), .A1(N18833), .B0(N18311), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11808 (.Y(N15794), .A0(N18672), .A1(N11207), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11809 (.Y(N15795), .A0(N18672), .A1(N8863), .B0(N18261), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11810 (.Y(N15796), .A0(N18677), .A1(N18739), .B0(N1044), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11811 (.Y(N15797), .A0(N18677), .A1(N14649), .B0(N11176), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11812 (.Y(N15798), .A0(N18677), .A1(N8867), .B0(N14658), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11813 (.Y(N15799), .A0(N18677), .A1(N11204), .B0(N4396), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11814 (.Y(N15800), .A0(N18677), .A1(N18400), .B0(N18259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11815 (.Y(N15801), .A0(N18677), .A1(N18407), .B0(N18725), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11816 (.Y(N15802), .A0(N18677), .A1(N18331), .B0(N18259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11818 (.Y(N15804), .A0(N18677), .A1(N18341), .B0(N18702), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11819 (.Y(N15805), .A0(N18677), .A1(N18341), .B0(N18583), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I12582 (.Y(N16832), .A(N18450), .B(N18911));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12589 (.Y(N16845), .A0(N18531), .A1(N18479), .B0(N18405), .B1(N18911));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I12601 (.Y(N16861), .A0(N18531), .A1(N18249), .B0(N18418), .B1(N18911));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12602 (.Y(N16862), .A0(N18531), .A1(N18430), .B0(N18400), .B1(N18911));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I12608 (.Y(N16869), .A(N18911), .B(N18249));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12612 (.Y(N16878), .A0(N18531), .A1(N18418), .B0(N18573), .B1(N18911));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I12613 (.Y(N16879), .A(N18531), .B(N18411));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12615 (.Y(N16882), .A0(N18531), .A1(N18400), .B0(N18405), .B1(N18911));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13383 (.Y(N17901), .A(N18466));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13390 (.Y(N17908), .A(N18411), .B(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13413 (.Y(N17948), .A0(N18531), .A1(N18221), .B0(N18460), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13416 (.Y(N17951), .A0(N18531), .A1(N18221), .B0(N18411), .B1(N18909));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13427 (.Y(N17969), .A0(N18677), .A1(N5555), .B0(N18241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13428 (.Y(N17970), .A0(N18672), .A1(N18739), .B0(N14658), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13429 (.Y(N17971), .A0(N18672), .A1(N18307), .B0(N6633), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13430 (.Y(N17972), .A0(N18672), .A1(N18725), .B0(N18231), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13431 (.Y(N17973), .A0(N18672), .A1(N18706), .B0(N18885), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13432 (.Y(N17974), .A0(N18672), .A1(N18259), .B0(N18407), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13433 (.Y(N17975), .A0(N18672), .A1(N18717), .B0(N18265), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13434 (.Y(N17976), .A0(N18672), .A1(N18583), .B0(N18253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13437 (.Y(N17982), .A0(N18672), .A1(N17901), .B0(N5593), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13438 (.Y(N17983), .A0(N18672), .A1(N18706), .B0(N16832), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13439 (.Y(N17984), .A0(N18672), .A1(N2141), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I13440 (.Y(N17985), .A0(N18672), .A1(N16861), .B0(N12316), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13441 (.Y(N17986), .A0(N18672), .A1(N14619), .B0(N18243), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13442 (.Y(N17987), .A(N18672), .B(N10146));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13443 (.Y(N17989), .A0(N18672), .A1(N8814), .B0(N18897), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13444 (.Y(N17990), .A0(N18672), .A1(N17908), .B0(N2176), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13445 (.Y(N17991), .A0(N18672), .A1(N1089), .B0(N16845), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13446 (.Y(N17992), .A0(N18672), .A1(N18307), .B0(N18229), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13447 (.Y(N17993), .A0(N18672), .A1(N11181), .B0(N18333), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13448 (.Y(N17994), .A0(N18672), .A1(N1068), .B0(N18406), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13449 (.Y(N17995), .A0(N18672), .A1(N18833), .B0(N18291), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13450 (.Y(N17996), .A0(N18897), .A1(N18672), .B0(N18335), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13451 (.Y(N17997), .A0(N18672), .A1(N18908), .B0(N18315), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13452 (.Y(N17998), .A(N18269), .B(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13455 (.Y(N18002), .A0(N18672), .A1(N18347), .B0(N14638), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13456 (.Y(N18003), .A0(N18672), .A1(N12363), .B0(N18601), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13457 (.Y(N18004), .A0(N18672), .A1(N1093), .B0(N16861), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13458 (.Y(N18005), .A0(N18672), .A1(N10134), .B0(N16862), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13459 (.Y(N18006), .A0(N18672), .A1(N7753), .B0(N4329), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13460 (.Y(N18007), .A0(N18672), .A1(N16878), .B0(N14649), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13461 (.Y(N18008), .A0(N18672), .A1(N18722), .B0(N18295), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13462 (.Y(N18009), .A0(N18672), .A1(N15724), .B0(N18301), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13463 (.Y(N18010), .A0(N18672), .A1(N11210), .B0(N8819), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13464 (.Y(N18011), .A0(N18672), .A1(N11176), .B0(N16869), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13465 (.Y(N18012), .A0(N18672), .A1(N3309), .B0(N4382), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13466 (.Y(N18013), .A0(N18672), .A1(N1045), .B0(N18261), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13467 (.Y(N18014), .A0(N18672), .A1(N17948), .B0(N18245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13468 (.Y(N18015), .A0(N18672), .A1(N18281), .B0(N16878), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13469 (.Y(N18016), .A0(N18672), .A1(N18295), .B0(N16879), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13470 (.Y(N18017), .A0(N18672), .A1(N17951), .B0(N12346), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13471 (.Y(N18018), .A0(N18672), .A1(N12363), .B0(N16882), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13472 (.Y(N18019), .A0(N18672), .A1(N18702), .B0(N3327), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13473 (.Y(N18020), .A(N18672), .B(N18327));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13474 (.Y(N18023), .A0(N18672), .A1(N18400), .B0(N18833), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13475 (.Y(N18024), .A0(N18672), .A1(N18406), .B0(N13459), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13476 (.Y(N18025), .A0(N18531), .A1(N18672), .B0(N18281), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13477 (.Y(N18026), .A(N18672), .B(N18596));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13481 (.Y(N18034), .A0(N18802), .A1(N17969), .B0(N15750), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13482 (.Y(N18035), .A0(N18802), .A1(N17970), .B0(N15751), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13483 (.Y(N18036), .A0(N18802), .A1(N17971), .B0(N15752), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13484 (.Y(N18037), .A0(N18802), .A1(N17972), .B0(N15753), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13485 (.Y(N18038), .A0(N18802), .A1(N17973), .B0(N15754), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13486 (.Y(N18039), .A0(N18802), .A1(N17974), .B0(N15755), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13487 (.Y(N18040), .A0(N18802), .A1(N17975), .B0(N15756), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13488 (.Y(N18041), .A0(N18802), .A1(N17976), .B0(N2203), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13491 (.Y(N18046), .A0(N18802), .A1(N17982), .B0(N15762), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13492 (.Y(N18047), .A0(N18802), .A1(N17983), .B0(N15763), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13493 (.Y(N18048), .A0(N18802), .A1(N17984), .B0(N15764), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13494 (.Y(N18049), .A0(N18802), .A1(N17985), .B0(N15765), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13495 (.Y(N18050), .A0(N18802), .A1(N17986), .B0(N15766), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13496 (.Y(N18051), .A0(N18802), .A1(N17987), .B0(N15767), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13497 (.Y(N18052), .A0(N18802), .A1(N17989), .B0(N15768), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13498 (.Y(N18053), .A0(N18802), .A1(N17990), .B0(N15769), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13499 (.Y(N18054), .A0(N18802), .A1(N17991), .B0(N15770), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13500 (.Y(N18055), .A0(N18802), .A1(N17992), .B0(N15771), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13501 (.Y(N18056), .A0(N18802), .A1(N17993), .B0(N15772), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13502 (.Y(N18057), .A0(N18802), .A1(N17994), .B0(N15773), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13503 (.Y(N18058), .A0(N18802), .A1(N17995), .B0(N15774), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13504 (.Y(N18059), .A0(N18802), .A1(N17996), .B0(N15775), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13505 (.Y(N18060), .A0(N18802), .A1(N17997), .B0(N15776), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13506 (.Y(N18061), .A0(N18802), .A1(N17998), .B0(N4473), .B1(N19085));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13507 (.Y(N18062), .A(N18802), .B(N4470));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13509 (.Y(N18067), .A0(N18802), .A1(N18002), .B0(N15783), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13510 (.Y(N18068), .A0(N18802), .A1(N18003), .B0(N15784), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13511 (.Y(N18069), .A0(N18802), .A1(N18004), .B0(N15785), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13512 (.Y(N18070), .A0(N18802), .A1(N18005), .B0(N15786), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13513 (.Y(N18071), .A0(N18802), .A1(N18006), .B0(N15787), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13514 (.Y(N18072), .A0(N18802), .A1(N18007), .B0(N15788), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13515 (.Y(N18073), .A0(N18802), .A1(N18008), .B0(N15789), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13516 (.Y(N18074), .A0(N18802), .A1(N18009), .B0(N15790), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13517 (.Y(N18075), .A0(N18802), .A1(N18010), .B0(N15791), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13518 (.Y(N18076), .A0(N18802), .A1(N18011), .B0(N15792), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13519 (.Y(N18077), .A0(N18802), .A1(N18012), .B0(N15793), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13520 (.Y(N18078), .A0(N18802), .A1(N18013), .B0(N15794), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13521 (.Y(N18079), .A0(N18802), .A1(N18014), .B0(N15795), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13522 (.Y(N18080), .A0(N18802), .A1(N18015), .B0(N15796), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13523 (.Y(N18081), .A0(N18802), .A1(N18016), .B0(N15797), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13524 (.Y(N18082), .A0(N18802), .A1(N18017), .B0(N15798), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13525 (.Y(N18083), .A0(N18802), .A1(N18018), .B0(N15799), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13526 (.Y(N18084), .A0(N18802), .A1(N18019), .B0(N15800), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13527 (.Y(N18085), .A0(N18802), .A1(N18020), .B0(N15801), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13528 (.Y(N18086), .A0(N18802), .A1(N18023), .B0(N15802), .B1(N19085));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13529 (.Y(N18087), .A0(N18802), .A1(N18024), .B0(N4436), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13530 (.Y(N18088), .A0(N18802), .A1(N18025), .B0(N15804), .B1(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13531 (.Y(N18089), .A0(N18802), .A1(N18026), .B0(N15805), .B1(N19086));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13532 (.Y(N18090), .A(N11243), .B(N19086));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13535 (.Y(N18094), .A0(N18865), .A1(N18034), .B0(N13538), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13536 (.Y(N18095), .A0(N18865), .A1(N18035), .B0(N13539), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13537 (.Y(N18096), .A0(N18865), .A1(N18036), .B0(N13540), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13538 (.Y(N18097), .A0(N18865), .A1(N18037), .B0(N13541), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13539 (.Y(N18098), .A0(N18865), .A1(N18038), .B0(N13542), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13540 (.Y(N18099), .A0(N18865), .A1(N18039), .B0(N13543), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13541 (.Y(N18100), .A0(N18865), .A1(N18040), .B0(N13544), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13542 (.Y(N18101), .A0(N18865), .A1(N18041), .B0(N13545), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13543 (.Y(N18102), .A0(N18865), .A1(N9022), .B0(N13546), .B1(N19111));
NOR2XL andori2bb1_A_I14593 (.Y(N19153), .A(N19085), .B(N2261));
NOR2XL andori2bb1_A_I14594 (.Y(N18103), .A(N19153), .B(N18865));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13545 (.Y(N18106), .A0(N18865), .A1(N18046), .B0(N13551), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13546 (.Y(N18107), .A0(N18865), .A1(N18047), .B0(N13552), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13547 (.Y(N18108), .A0(N18865), .A1(N18048), .B0(N13553), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13548 (.Y(N18109), .A0(N18865), .A1(N18049), .B0(N13554), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13549 (.Y(N18110), .A0(N18865), .A1(N18050), .B0(N13555), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13550 (.Y(N18111), .A0(N18865), .A1(N18051), .B0(N13556), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13551 (.Y(N18112), .A0(N18865), .A1(N18052), .B0(N13557), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13552 (.Y(N18113), .A0(N18865), .A1(N18053), .B0(N13558), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13553 (.Y(N18114), .A0(N18865), .A1(N18054), .B0(N13559), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13554 (.Y(N18115), .A0(N18865), .A1(N18055), .B0(N13560), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13555 (.Y(N18116), .A0(N18865), .A1(N18056), .B0(N13561), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13556 (.Y(N18117), .A0(N18865), .A1(N18057), .B0(N13562), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13557 (.Y(N18118), .A0(N18865), .A1(N18058), .B0(N13563), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13558 (.Y(N18119), .A0(N18865), .A1(N18059), .B0(N13564), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13559 (.Y(N18120), .A0(N18865), .A1(N18060), .B0(N13565), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13560 (.Y(N18121), .A0(N18865), .A1(N18061), .B0(N13566), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13561 (.Y(N18122), .A0(N18865), .A1(N18062), .B0(N13567), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13563 (.Y(N18125), .A0(N18865), .A1(N18067), .B0(N13572), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13564 (.Y(N18126), .A0(N18865), .A1(N18068), .B0(N13573), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13565 (.Y(N18127), .A0(N18865), .A1(N18069), .B0(N13574), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13566 (.Y(N18128), .A0(N18865), .A1(N18070), .B0(N13575), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13567 (.Y(N18129), .A0(N18865), .A1(N18071), .B0(N13576), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13568 (.Y(N18130), .A0(N18865), .A1(N18072), .B0(N13577), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13569 (.Y(N18131), .A0(N18865), .A1(N18073), .B0(N13578), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13570 (.Y(N18132), .A0(N18865), .A1(N18074), .B0(N13579), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13571 (.Y(N18133), .A0(N18865), .A1(N18075), .B0(N13580), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13572 (.Y(N18134), .A0(N18865), .A1(N18076), .B0(N13581), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13573 (.Y(N18135), .A0(N18865), .A1(N18077), .B0(N13582), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13574 (.Y(N18136), .A0(N18865), .A1(N18078), .B0(N13583), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13575 (.Y(N18137), .A0(N18865), .A1(N18079), .B0(N13584), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13576 (.Y(N18138), .A0(N18865), .A1(N18080), .B0(N13585), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13577 (.Y(N18139), .A0(N18865), .A1(N18081), .B0(N13586), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13578 (.Y(N18140), .A0(N18865), .A1(N18082), .B0(N13587), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13579 (.Y(N18141), .A0(N18865), .A1(N18083), .B0(N13588), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13580 (.Y(N18142), .A0(N18865), .A1(N18084), .B0(N13589), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13581 (.Y(N18143), .A0(N18865), .A1(N18085), .B0(N13590), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13582 (.Y(N18144), .A0(N18865), .A1(N18086), .B0(N13591), .B1(N19111));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13583 (.Y(N18145), .A0(N18865), .A1(N18087), .B0(N13592), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13584 (.Y(N18146), .A0(N18865), .A1(N18088), .B0(N13593), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13585 (.Y(N18147), .A0(N18865), .A1(N18089), .B0(N13594), .B1(N19112));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13586 (.Y(N18148), .A0(N18865), .A1(N18090), .B0(N8968), .B1(N19112));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14209 (.Y(N18880), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13589 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[0]), .A0(N18880), .A1(N18094), .B0(N9028), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13590 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[1]), .A0(N18880), .A1(N18095), .B0(N9029), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13591 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[2]), .A0(N18880), .A1(N18096), .B0(N9030), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13592 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[3]), .A0(N18880), .A1(N18097), .B0(N9031), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13593 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[4]), .A0(N18880), .A1(N18098), .B0(N9032), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13594 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[5]), .A0(N18880), .A1(N18099), .B0(N9033), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13595 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[6]), .A0(N18880), .A1(N18100), .B0(N9034), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13596 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[7]), .A0(N18880), .A1(N18101), .B0(N9036), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13597 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[8]), .A0(N18880), .A1(N18102), .B0(N9039), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13598 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[9]), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]), .B(N18103));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13599 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[10]), .A0(N18880), .A1(N18106), .B0(N9042), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13600 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[11]), .A0(N18880), .A1(N18107), .B0(N9043), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13601 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[12]), .A0(N18880), .A1(N18108), .B0(N9044), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13602 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[13]), .A0(N18880), .A1(N18109), .B0(N9045), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13603 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[14]), .A0(N18880), .A1(N18110), .B0(N9046), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13604 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[15]), .A0(N18880), .A1(N18111), .B0(N9047), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13605 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[16]), .A0(N18880), .A1(N18112), .B0(N9048), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13606 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[17]), .A0(N18880), .A1(N18113), .B0(N9049), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13607 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[18]), .A0(N18880), .A1(N18114), .B0(N9050), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13608 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[19]), .A0(N18880), .A1(N18115), .B0(N9051), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13609 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[20]), .A0(N18880), .A1(N18116), .B0(N9052), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13610 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[21]), .A0(N18880), .A1(N18117), .B0(N9053), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13611 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[22]), .A0(N18880), .A1(N18118), .B0(N9054), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13612 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[23]), .A0(N18880), .A1(N18119), .B0(N9055), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13613 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[24]), .A0(N18880), .A1(N18120), .B0(N9056), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13614 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[25]), .A0(N18880), .A1(N18121), .B0(N9057), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13615 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[26]), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]), .B(N18122));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I14523 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[27]), .A0N(N13569), .A1N(N19112), .B0(N18880));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13617 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[28]), .A0(N18880), .A1(N18125), .B0(N9063), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13618 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[29]), .A0(N18880), .A1(N18126), .B0(N9064), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13619 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[30]), .A0(N18880), .A1(N18127), .B0(N9065), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13620 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[31]), .A0(N18880), .A1(N18128), .B0(N9066), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13621 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[32]), .A0(N18880), .A1(N18129), .B0(N9067), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13622 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[33]), .A0(N18880), .A1(N18130), .B0(N9068), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13623 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[34]), .A0(N18880), .A1(N18131), .B0(N9069), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13624 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[35]), .A0(N18880), .A1(N18132), .B0(N9070), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13625 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[36]), .A0(N18880), .A1(N18133), .B0(N9071), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13626 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[37]), .A0(N18880), .A1(N18134), .B0(N9072), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13627 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[38]), .A0(N18880), .A1(N18135), .B0(N9073), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13628 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[39]), .A0(N18880), .A1(N18136), .B0(N9074), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13629 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[40]), .A0(N18880), .A1(N18137), .B0(N9075), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13630 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[41]), .A0(N18880), .A1(N18138), .B0(N9076), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13631 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[42]), .A0(N18880), .A1(N18139), .B0(N9077), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13632 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[43]), .A0(N18880), .A1(N18140), .B0(N9078), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13633 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[44]), .A0(N18880), .A1(N18141), .B0(N9079), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13634 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[45]), .A0(N18880), .A1(N18142), .B0(N9080), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13635 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[46]), .A0(N18880), .A1(N18143), .B0(N9081), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13636 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[47]), .A0(N18880), .A1(N18144), .B0(N9082), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13637 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[48]), .A0(N18880), .A1(N18145), .B0(N9083), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13638 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[49]), .A0(N18880), .A1(N18146), .B0(N9084), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13639 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[50]), .A0(N18880), .A1(N18147), .B0(N9085), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13640 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[51]), .A0(N18880), .A1(N18148), .B0(N9086), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL andori2bb1_A_I14595 (.Y(N19160), .A(N18865), .B(N8972));
NOR2XL andori2bb1_A_I14596 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[52]), .A(N19160), .B(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
endmodule

module cynw_cm_float_rcp_inst_cellmath__62_0_bdw1471647203_bdw (
	inst_cellmath__62_0_out0,
	inst_cellmath__62_0_out1,
	inst_cellmath__62_0_in0,
	inst_cellmath__62_0_in1
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__62_0_out0,
	inst_cellmath__62_0_out1;
input [9:0] inst_cellmath__62_0_in0;
input [24:13] inst_cellmath__62_0_in1;
wire N313,N315,N317,N319,N321,N323,N325 
	,N327,N329,N331,N346,N348,N350,N352,N354 
	,N356,N358,N360,N362,N364,N366,N381,N383 
	,N385,N387,N389,N391,N393,N395,N397,N399 
	,N401,N414,N416,N418,N420,N422,N424,N426 
	,N428,N430,N432,N434,N436,N449,N451,N453 
	,N455,N457,N459,N461,N463,N465,N467,N469 
	,N471,N484,N486,N488,N490,N492,N494,N496 
	,N498,N500,N502,N504,N506,N519,N521,N523 
	,N525,N527,N529,N531,N533,N535,N537,N539 
	,N541,N554,N556,N558,N560,N562,N564,N566 
	,N568,N570,N572,N574,N576,N589,N591,N593 
	,N595,N597,N599,N601,N603,N605,N607,N609 
	,N611,N624,N626,N628,N630,N632,N634,N636 
	,N638,N640,N642,N644,N650,N652,N654,N655 
	,N656,N658,N661,N662,N663,N664,N665,N666 
	,N669,N670,N671,N672,N673,N674,N675,N676 
	,N679,N680,N681,N682,N683,N684,N685,N686 
	,N687,N688,N691,N692,N693,N694,N695,N696 
	,N697,N698,N699,N700,N701,N702,N705,N706 
	,N707,N708,N709,N710,N711,N712,N713,N714 
	,N715,N716,N717,N718,N721,N722,N723,N724 
	,N725,N726,N727,N728,N729,N730,N731,N732 
	,N733,N734,N737,N738,N739,N740,N741,N742 
	,N743,N744,N745,N746,N747,N748,N749,N750 
	,N753,N754,N755,N756,N757,N758,N759,N760 
	,N761,N762,N763,N764,N765,N766,N769,N770 
	,N771,N772,N773,N774,N775,N776,N777,N778 
	,N779,N780,N783,N784,N785,N786,N787,N788 
	,N789,N790,N791,N792,N795,N796,N797,N798 
	,N799,N800,N801,N802,N805,N806,N807,N808 
	,N809,N810,N813,N814,N815,N816,N819,N820 
	,N825,N826,N827,N828,N829,N830,N831,N832 
	,N833,N834,N835,N836,N837,N838,N839,N840 
	,N841,N842,N843,N844,N845,N846;
INVX1 inst_cellmath__62_0_I303 (.Y(N825), .A(inst_cellmath__62_0_in1[13]));
INVXL inst_cellmath__62_0_I304 (.Y(N826), .A(inst_cellmath__62_0_in1[14]));
INVXL inst_cellmath__62_0_I305 (.Y(N827), .A(inst_cellmath__62_0_in1[15]));
INVX1 inst_cellmath__62_0_I306 (.Y(N828), .A(inst_cellmath__62_0_in1[16]));
INVX2 inst_cellmath__62_0_I307 (.Y(N829), .A(inst_cellmath__62_0_in1[17]));
INVXL inst_cellmath__62_0_I308 (.Y(N830), .A(inst_cellmath__62_0_in1[18]));
INVX3 inst_cellmath__62_0_I309 (.Y(N831), .A(inst_cellmath__62_0_in1[19]));
INVXL inst_cellmath__62_0_I310 (.Y(N832), .A(inst_cellmath__62_0_in1[20]));
INVX1 inst_cellmath__62_0_I311 (.Y(N833), .A(inst_cellmath__62_0_in1[21]));
INVX1 inst_cellmath__62_0_I312 (.Y(N834), .A(inst_cellmath__62_0_in1[22]));
INVXL inst_cellmath__62_0_I313 (.Y(N835), .A(inst_cellmath__62_0_in1[23]));
INVX1 inst_cellmath__62_0_I314 (.Y(N836), .A(inst_cellmath__62_0_in1[24]));
INVXL inst_cellmath__62_0_I315 (.Y(N837), .A(inst_cellmath__62_0_in0[0]));
NOR2XL inst_cellmath__62_0_I49 (.Y(inst_cellmath__62_0_out1[4]), .A(N837), .B(N825));
NOR2XL inst_cellmath__62_0_I50 (.Y(inst_cellmath__62_0_out1[5]), .A(N837), .B(N826));
NOR2XL inst_cellmath__62_0_I51 (.Y(N313), .A(N837), .B(N827));
NOR2XL inst_cellmath__62_0_I52 (.Y(N315), .A(N837), .B(N828));
NOR2XL inst_cellmath__62_0_I53 (.Y(N317), .A(N837), .B(N829));
NOR2XL inst_cellmath__62_0_I54 (.Y(N319), .A(N837), .B(N830));
NOR2XL inst_cellmath__62_0_I55 (.Y(N321), .A(N837), .B(N831));
NOR2XL inst_cellmath__62_0_I56 (.Y(N323), .A(N837), .B(N832));
NOR2XL inst_cellmath__62_0_I57 (.Y(N325), .A(N837), .B(N833));
NOR2XL inst_cellmath__62_0_I58 (.Y(N327), .A(N837), .B(N834));
NOR2XL inst_cellmath__62_0_I59 (.Y(N329), .A(N837), .B(N835));
NOR2XL inst_cellmath__62_0_I60 (.Y(N331), .A(N837), .B(N836));
INVXL inst_cellmath__62_0_I316 (.Y(N838), .A(inst_cellmath__62_0_in0[1]));
NOR2XL inst_cellmath__62_0_I66 (.Y(inst_cellmath__62_0_out0[5]), .A(N838), .B(N825));
NOR2XL inst_cellmath__62_0_I67 (.Y(N346), .A(N838), .B(N826));
NOR2XL inst_cellmath__62_0_I68 (.Y(N348), .A(N838), .B(N827));
NOR2XL inst_cellmath__62_0_I69 (.Y(N350), .A(N838), .B(N828));
NOR2XL inst_cellmath__62_0_I70 (.Y(N352), .A(N838), .B(N829));
NOR2XL inst_cellmath__62_0_I71 (.Y(N354), .A(N838), .B(N830));
NOR2XL inst_cellmath__62_0_I72 (.Y(N356), .A(N838), .B(N831));
NOR2XL inst_cellmath__62_0_I73 (.Y(N358), .A(N838), .B(N832));
NOR2XL inst_cellmath__62_0_I74 (.Y(N360), .A(N838), .B(N833));
NOR2XL inst_cellmath__62_0_I75 (.Y(N362), .A(N838), .B(N834));
NOR2XL inst_cellmath__62_0_I76 (.Y(N364), .A(N838), .B(N835));
NOR2XL inst_cellmath__62_0_I77 (.Y(N366), .A(N838), .B(N836));
INVXL inst_cellmath__62_0_I317 (.Y(N839), .A(inst_cellmath__62_0_in0[2]));
NOR2XL inst_cellmath__62_0_I83 (.Y(inst_cellmath__62_0_out1[6]), .A(N839), .B(N825));
NOR2XL inst_cellmath__62_0_I84 (.Y(N381), .A(N839), .B(N826));
NOR2XL inst_cellmath__62_0_I85 (.Y(N383), .A(N839), .B(N827));
NOR2XL inst_cellmath__62_0_I86 (.Y(N385), .A(N839), .B(N828));
NOR2XL inst_cellmath__62_0_I87 (.Y(N387), .A(N839), .B(N829));
NOR2XL inst_cellmath__62_0_I88 (.Y(N389), .A(N839), .B(N830));
NOR2XL inst_cellmath__62_0_I89 (.Y(N391), .A(N839), .B(N831));
NOR2XL inst_cellmath__62_0_I90 (.Y(N393), .A(N839), .B(N832));
NOR2XL inst_cellmath__62_0_I91 (.Y(N395), .A(N839), .B(N833));
NOR2XL inst_cellmath__62_0_I92 (.Y(N397), .A(N839), .B(N834));
NOR2XL inst_cellmath__62_0_I93 (.Y(N399), .A(N839), .B(N835));
NOR2XL inst_cellmath__62_0_I94 (.Y(N401), .A(N839), .B(N836));
INVXL inst_cellmath__62_0_I318 (.Y(N840), .A(inst_cellmath__62_0_in0[3]));
NOR2XL inst_cellmath__62_0_I100 (.Y(N414), .A(N840), .B(N825));
NOR2XL inst_cellmath__62_0_I101 (.Y(N416), .A(N840), .B(N826));
NOR2XL inst_cellmath__62_0_I102 (.Y(N418), .A(N840), .B(N827));
NOR2XL inst_cellmath__62_0_I103 (.Y(N420), .A(N840), .B(N828));
NOR2XL inst_cellmath__62_0_I104 (.Y(N422), .A(N840), .B(N829));
NOR2XL inst_cellmath__62_0_I105 (.Y(N424), .A(N840), .B(N830));
NOR2XL inst_cellmath__62_0_I106 (.Y(N426), .A(N840), .B(N831));
NOR2XL inst_cellmath__62_0_I107 (.Y(N428), .A(N840), .B(N832));
NOR2XL inst_cellmath__62_0_I108 (.Y(N430), .A(N840), .B(N833));
NOR2XL inst_cellmath__62_0_I109 (.Y(N432), .A(N840), .B(N834));
NOR2XL inst_cellmath__62_0_I110 (.Y(N434), .A(N840), .B(N835));
NOR2XL inst_cellmath__62_0_I111 (.Y(N436), .A(N840), .B(N836));
INVXL inst_cellmath__62_0_I319 (.Y(N841), .A(inst_cellmath__62_0_in0[4]));
NOR2XL inst_cellmath__62_0_I117 (.Y(N449), .A(N841), .B(N825));
NOR2XL inst_cellmath__62_0_I118 (.Y(N451), .A(N841), .B(N826));
NOR2XL inst_cellmath__62_0_I119 (.Y(N453), .A(N841), .B(N827));
NOR2XL inst_cellmath__62_0_I120 (.Y(N455), .A(N841), .B(N828));
NOR2XL inst_cellmath__62_0_I121 (.Y(N457), .A(N841), .B(N829));
NOR2XL inst_cellmath__62_0_I122 (.Y(N459), .A(N841), .B(N830));
NOR2X1 inst_cellmath__62_0_I123 (.Y(N461), .A(N841), .B(N831));
NOR2XL inst_cellmath__62_0_I124 (.Y(N463), .A(N841), .B(N832));
NOR2XL inst_cellmath__62_0_I125 (.Y(N465), .A(N841), .B(N833));
NOR2XL inst_cellmath__62_0_I126 (.Y(N467), .A(N841), .B(N834));
NOR2XL inst_cellmath__62_0_I127 (.Y(N469), .A(N841), .B(N835));
NOR2XL inst_cellmath__62_0_I128 (.Y(N471), .A(N841), .B(N836));
INVXL inst_cellmath__62_0_I320 (.Y(N842), .A(inst_cellmath__62_0_in0[5]));
NOR2XL inst_cellmath__62_0_I134 (.Y(N484), .A(N842), .B(N825));
NOR2XL inst_cellmath__62_0_I135 (.Y(N486), .A(N842), .B(N826));
NOR2XL inst_cellmath__62_0_I136 (.Y(N488), .A(N842), .B(N827));
NOR2XL inst_cellmath__62_0_I137 (.Y(N490), .A(N842), .B(N828));
NOR2XL inst_cellmath__62_0_I138 (.Y(N492), .A(N842), .B(N829));
NOR2XL inst_cellmath__62_0_I139 (.Y(N494), .A(N842), .B(N830));
NOR2XL inst_cellmath__62_0_I140 (.Y(N496), .A(N842), .B(N831));
NOR2XL inst_cellmath__62_0_I141 (.Y(N498), .A(N842), .B(N832));
NOR2XL inst_cellmath__62_0_I142 (.Y(N500), .A(N842), .B(N833));
NOR2XL inst_cellmath__62_0_I143 (.Y(N502), .A(N842), .B(N834));
NOR2XL inst_cellmath__62_0_I144 (.Y(N504), .A(N842), .B(N835));
NOR2XL inst_cellmath__62_0_I145 (.Y(N506), .A(N842), .B(N836));
INVXL inst_cellmath__62_0_I321 (.Y(N843), .A(inst_cellmath__62_0_in0[6]));
NOR2XL inst_cellmath__62_0_I151 (.Y(N519), .A(N843), .B(N825));
NOR2XL inst_cellmath__62_0_I152 (.Y(N521), .A(N843), .B(N826));
NOR2XL inst_cellmath__62_0_I153 (.Y(N523), .A(N843), .B(N827));
NOR2XL inst_cellmath__62_0_I154 (.Y(N525), .A(N843), .B(N828));
NOR2XL inst_cellmath__62_0_I155 (.Y(N527), .A(N843), .B(N829));
NOR2XL inst_cellmath__62_0_I156 (.Y(N529), .A(N843), .B(N830));
NOR2X1 inst_cellmath__62_0_I157 (.Y(N531), .A(N843), .B(N831));
NOR2XL inst_cellmath__62_0_I158 (.Y(N533), .A(N843), .B(N832));
NOR2XL inst_cellmath__62_0_I159 (.Y(N535), .A(N843), .B(N833));
NOR2XL inst_cellmath__62_0_I160 (.Y(N537), .A(N843), .B(N834));
NOR2XL inst_cellmath__62_0_I161 (.Y(N539), .A(N843), .B(N835));
NOR2XL inst_cellmath__62_0_I162 (.Y(N541), .A(N843), .B(N836));
INVXL inst_cellmath__62_0_I322 (.Y(N844), .A(inst_cellmath__62_0_in0[7]));
NOR2XL inst_cellmath__62_0_I168 (.Y(N554), .A(N844), .B(N825));
NOR2XL inst_cellmath__62_0_I169 (.Y(N556), .A(N844), .B(N826));
NOR2XL inst_cellmath__62_0_I170 (.Y(N558), .A(N844), .B(N827));
NOR2XL inst_cellmath__62_0_I171 (.Y(N560), .A(N844), .B(N828));
NOR2XL inst_cellmath__62_0_I172 (.Y(N562), .A(N844), .B(N829));
NOR2XL inst_cellmath__62_0_I173 (.Y(N564), .A(N844), .B(N830));
NOR2XL inst_cellmath__62_0_I174 (.Y(N566), .A(N844), .B(N831));
NOR2XL inst_cellmath__62_0_I175 (.Y(N568), .A(N844), .B(N832));
NOR2XL inst_cellmath__62_0_I176 (.Y(N570), .A(N844), .B(N833));
NOR2XL inst_cellmath__62_0_I177 (.Y(N572), .A(N844), .B(N834));
NOR2XL inst_cellmath__62_0_I178 (.Y(N574), .A(N844), .B(N835));
NOR2XL inst_cellmath__62_0_I179 (.Y(N576), .A(N844), .B(N836));
INVXL inst_cellmath__62_0_I323 (.Y(N845), .A(inst_cellmath__62_0_in0[8]));
NOR2XL inst_cellmath__62_0_I185 (.Y(N589), .A(N845), .B(N825));
NOR2XL inst_cellmath__62_0_I186 (.Y(N591), .A(N845), .B(N826));
NOR2XL inst_cellmath__62_0_I187 (.Y(N593), .A(N845), .B(N827));
NOR2XL inst_cellmath__62_0_I188 (.Y(N595), .A(N845), .B(N828));
NOR2XL inst_cellmath__62_0_I189 (.Y(N597), .A(N845), .B(N829));
NOR2XL inst_cellmath__62_0_I190 (.Y(N599), .A(N845), .B(N830));
NOR2XL inst_cellmath__62_0_I191 (.Y(N601), .A(N845), .B(N831));
NOR2XL inst_cellmath__62_0_I192 (.Y(N603), .A(N845), .B(N832));
NOR2XL inst_cellmath__62_0_I193 (.Y(N605), .A(N845), .B(N833));
NOR2XL inst_cellmath__62_0_I194 (.Y(N607), .A(N845), .B(N834));
NOR2XL inst_cellmath__62_0_I195 (.Y(N609), .A(N845), .B(N835));
NOR2XL inst_cellmath__62_0_I196 (.Y(N611), .A(N845), .B(N836));
INVXL inst_cellmath__62_0_I324 (.Y(N846), .A(inst_cellmath__62_0_in0[9]));
NOR2XL inst_cellmath__62_0_I202 (.Y(N624), .A(N846), .B(N825));
NOR2XL inst_cellmath__62_0_I203 (.Y(N626), .A(N846), .B(N826));
NOR2XL inst_cellmath__62_0_I204 (.Y(N628), .A(N846), .B(N827));
NOR2XL inst_cellmath__62_0_I205 (.Y(N630), .A(N846), .B(N828));
NOR2XL inst_cellmath__62_0_I206 (.Y(N632), .A(N846), .B(N829));
NOR2XL inst_cellmath__62_0_I207 (.Y(N634), .A(N846), .B(N830));
NOR2XL inst_cellmath__62_0_I208 (.Y(N636), .A(N846), .B(N831));
NOR2XL inst_cellmath__62_0_I209 (.Y(N638), .A(N846), .B(N832));
NOR2XL inst_cellmath__62_0_I210 (.Y(N640), .A(N846), .B(N833));
NOR2XL inst_cellmath__62_0_I211 (.Y(N642), .A(N846), .B(N834));
NOR2XL inst_cellmath__62_0_I212 (.Y(N644), .A(N846), .B(N835));
NOR2XL inst_cellmath__62_0_I213 (.Y(inst_cellmath__62_0_out1[24]), .A(N846), .B(N836));
ADDHX1 inst_cellmath__62_0_I215 (.CO(N650), .S(inst_cellmath__62_0_out0[6]), .A(N346), .B(N313));
ADDHX1 inst_cellmath__62_0_I216 (.CO(N652), .S(inst_cellmath__62_0_out1[7]), .A(N315), .B(N414));
ADDFX1 inst_cellmath__62_0_I217 (.CO(N654), .S(inst_cellmath__62_0_out0[7]), .A(N348), .B(N381), .CI(N650));
ADDHX1 inst_cellmath__62_0_I218 (.CO(N656), .S(N655), .A(N350), .B(N317));
ADDFX1 inst_cellmath__62_0_I219 (.CO(N658), .S(inst_cellmath__62_0_out1[8]), .A(N449), .B(N416), .CI(N383));
ADDFX1 inst_cellmath__62_0_I220 (.CO(inst_cellmath__62_0_out1[9]), .S(inst_cellmath__62_0_out0[8]), .A(N655), .B(N652), .CI(N654));
ADDHX1 inst_cellmath__62_0_I221 (.CO(N662), .S(N661), .A(N385), .B(N352));
ADDFX1 inst_cellmath__62_0_I222 (.CO(N664), .S(N663), .A(N484), .B(N451), .CI(N319));
ADDFX1 inst_cellmath__62_0_I223 (.CO(N666), .S(N665), .A(N656), .B(N418), .CI(N661));
ADDFX1 inst_cellmath__62_0_I224 (.CO(inst_cellmath__62_0_out1[10]), .S(inst_cellmath__62_0_out0[9]), .A(N663), .B(N658), .CI(N665));
ADDHX1 inst_cellmath__62_0_I225 (.CO(N670), .S(N669), .A(N420), .B(N387));
ADDFX1 inst_cellmath__62_0_I226 (.CO(N672), .S(N671), .A(N519), .B(N486), .CI(N354));
ADDFX1 inst_cellmath__62_0_I227 (.CO(N674), .S(N673), .A(N321), .B(N453), .CI(N662));
ADDFX1 inst_cellmath__62_0_I228 (.CO(N676), .S(N675), .A(N664), .B(N669), .CI(N671));
ADDFX1 inst_cellmath__62_0_I229 (.CO(inst_cellmath__62_0_out1[11]), .S(inst_cellmath__62_0_out0[10]), .A(N673), .B(N666), .CI(N675));
ADDHX1 inst_cellmath__62_0_I230 (.CO(N680), .S(N679), .A(N455), .B(N422));
ADDFX1 inst_cellmath__62_0_I231 (.CO(N682), .S(N681), .A(N554), .B(N521), .CI(N389));
ADDFX1 inst_cellmath__62_0_I232 (.CO(N684), .S(N683), .A(N356), .B(N488), .CI(N323));
ADDFX1 inst_cellmath__62_0_I233 (.CO(N686), .S(N685), .A(N679), .B(N670), .CI(N672));
ADDFX1 inst_cellmath__62_0_I234 (.CO(N688), .S(N687), .A(N681), .B(N674), .CI(N683));
ADDFX1 inst_cellmath__62_0_I235 (.CO(inst_cellmath__62_0_out1[12]), .S(inst_cellmath__62_0_out0[11]), .A(N685), .B(N676), .CI(N687));
ADDHX1 inst_cellmath__62_0_I236 (.CO(N692), .S(N691), .A(N490), .B(N457));
ADDFX1 inst_cellmath__62_0_I237 (.CO(N694), .S(N693), .A(N589), .B(N556), .CI(N424));
ADDFX1 inst_cellmath__62_0_I238 (.CO(N696), .S(N695), .A(N391), .B(N523), .CI(N358));
ADDFX1 inst_cellmath__62_0_I239 (.CO(N698), .S(N697), .A(N325), .B(N680), .CI(N691));
ADDFX1 inst_cellmath__62_0_I240 (.CO(N700), .S(N699), .A(N684), .B(N682), .CI(N693));
ADDFX1 inst_cellmath__62_0_I241 (.CO(N702), .S(N701), .A(N686), .B(N695), .CI(N697));
ADDFX1 inst_cellmath__62_0_I242 (.CO(inst_cellmath__62_0_out1[13]), .S(inst_cellmath__62_0_out0[12]), .A(N699), .B(N688), .CI(N701));
ADDHX1 inst_cellmath__62_0_I243 (.CO(N706), .S(N705), .A(N525), .B(N492));
ADDFX1 inst_cellmath__62_0_I244 (.CO(N708), .S(N707), .A(N624), .B(N591), .CI(N459));
ADDFX1 inst_cellmath__62_0_I245 (.CO(N710), .S(N709), .A(N426), .B(N558), .CI(N393));
ADDFX1 inst_cellmath__62_0_I246 (.CO(N712), .S(N711), .A(N692), .B(N327), .CI(N360));
ADDFX1 inst_cellmath__62_0_I247 (.CO(N714), .S(N713), .A(N694), .B(N705), .CI(N696));
ADDFX1 inst_cellmath__62_0_I248 (.CO(N716), .S(N715), .A(N698), .B(N707), .CI(N709));
ADDFX1 inst_cellmath__62_0_I249 (.CO(N718), .S(N717), .A(N700), .B(N711), .CI(N713));
ADDFX1 inst_cellmath__62_0_I250 (.CO(inst_cellmath__62_0_out1[14]), .S(inst_cellmath__62_0_out0[13]), .A(N715), .B(N702), .CI(N717));
ADDFX1 inst_cellmath__62_0_I251 (.CO(N722), .S(N721), .A(N626), .B(N560), .CI(N494));
ADDFX1 inst_cellmath__62_0_I252 (.CO(N724), .S(N723), .A(N461), .B(N527), .CI(N593));
ADDFX1 inst_cellmath__62_0_I253 (.CO(N726), .S(N725), .A(N362), .B(N428), .CI(N329));
ADDFX1 inst_cellmath__62_0_I254 (.CO(N728), .S(N727), .A(N395), .B(N706), .CI(N708));
ADDFX1 inst_cellmath__62_0_I255 (.CO(N730), .S(N729), .A(N721), .B(N710), .CI(N712));
ADDFX1 inst_cellmath__62_0_I256 (.CO(N732), .S(N731), .A(N725), .B(N723), .CI(N714));
ADDFX1 inst_cellmath__62_0_I257 (.CO(N734), .S(N733), .A(N716), .B(N727), .CI(N729));
ADDFX1 inst_cellmath__62_0_I258 (.CO(inst_cellmath__62_0_out1[15]), .S(inst_cellmath__62_0_out0[14]), .A(N731), .B(N718), .CI(N733));
ADDFX1 inst_cellmath__62_0_I259 (.CO(N738), .S(N737), .A(N529), .B(N595), .CI(N562));
ADDFX1 inst_cellmath__62_0_I260 (.CO(N740), .S(N739), .A(N496), .B(N628), .CI(N463));
ADDFX1 inst_cellmath__62_0_I261 (.CO(N742), .S(N741), .A(N397), .B(N331), .CI(N430));
ADDFX1 inst_cellmath__62_0_I262 (.CO(N744), .S(N743), .A(N722), .B(N364), .CI(N724));
ADDFX1 inst_cellmath__62_0_I263 (.CO(N746), .S(N745), .A(N726), .B(N737), .CI(N739));
ADDFX1 inst_cellmath__62_0_I264 (.CO(N748), .S(N747), .A(N741), .B(N728), .CI(N730));
ADDFX1 inst_cellmath__62_0_I265 (.CO(N750), .S(N749), .A(N732), .B(N743), .CI(N745));
ADDFX1 inst_cellmath__62_0_I266 (.CO(inst_cellmath__62_0_out1[16]), .S(inst_cellmath__62_0_out0[15]), .A(N747), .B(N734), .CI(N749));
ADDHX1 inst_cellmath__62_0_I267 (.CO(N754), .S(N753), .A(N630), .B(N597));
ADDFX1 inst_cellmath__62_0_I268 (.CO(N756), .S(N755), .A(N531), .B(N564), .CI(N498));
ADDFX1 inst_cellmath__62_0_I269 (.CO(N758), .S(N757), .A(N432), .B(N366), .CI(N465));
ADDFX1 inst_cellmath__62_0_I270 (.CO(N760), .S(N759), .A(N753), .B(N399), .CI(N738));
ADDFX1 inst_cellmath__62_0_I271 (.CO(N762), .S(N761), .A(N742), .B(N740), .CI(N755));
ADDFX1 inst_cellmath__62_0_I272 (.CO(N764), .S(N763), .A(N744), .B(N757), .CI(N759));
ADDFX1 inst_cellmath__62_0_I273 (.CO(N766), .S(N765), .A(N761), .B(N746), .CI(N748));
ADDFX1 inst_cellmath__62_0_I274 (.CO(inst_cellmath__62_0_out1[17]), .S(inst_cellmath__62_0_out0[16]), .A(N750), .B(N763), .CI(N765));
ADDFX1 inst_cellmath__62_0_I275 (.CO(N770), .S(N769), .A(N632), .B(N599), .CI(N566));
ADDFX1 inst_cellmath__62_0_I276 (.CO(N772), .S(N771), .A(N401), .B(N533), .CI(N467));
ADDFX1 inst_cellmath__62_0_I277 (.CO(N774), .S(N773), .A(N500), .B(N754), .CI(N434));
ADDFX1 inst_cellmath__62_0_I278 (.CO(N776), .S(N775), .A(N758), .B(N756), .CI(N769));
ADDFX1 inst_cellmath__62_0_I279 (.CO(N778), .S(N777), .A(N771), .B(N760), .CI(N773));
ADDFXL inst_cellmath__62_0_I280 (.CO(N780), .S(N779), .A(N775), .B(N762), .CI(N764));
ADDFXL inst_cellmath__62_0_I281 (.CO(inst_cellmath__62_0_out1[18]), .S(inst_cellmath__62_0_out0[17]), .A(N766), .B(N777), .CI(N779));
ADDFX1 inst_cellmath__62_0_I282 (.CO(N784), .S(N783), .A(N601), .B(N634), .CI(N568));
ADDFX1 inst_cellmath__62_0_I283 (.CO(N786), .S(N785), .A(N502), .B(N436), .CI(N535));
ADDFX1 inst_cellmath__62_0_I284 (.CO(N788), .S(N787), .A(N770), .B(N469), .CI(N772));
ADDFX1 inst_cellmath__62_0_I285 (.CO(N790), .S(N789), .A(N783), .B(N774), .CI(N785));
ADDFX1 inst_cellmath__62_0_I286 (.CO(N792), .S(N791), .A(N787), .B(N776), .CI(N778));
ADDFXL inst_cellmath__62_0_I287 (.CO(inst_cellmath__62_0_out1[19]), .S(inst_cellmath__62_0_out0[18]), .A(N780), .B(N789), .CI(N791));
ADDFX1 inst_cellmath__62_0_I288 (.CO(N796), .S(N795), .A(N603), .B(N636), .CI(N471));
ADDFX1 inst_cellmath__62_0_I289 (.CO(N798), .S(N797), .A(N570), .B(N537), .CI(N504));
ADDFX1 inst_cellmath__62_0_I290 (.CO(N800), .S(N799), .A(N786), .B(N784), .CI(N795));
ADDFXL inst_cellmath__62_0_I291 (.CO(N802), .S(N801), .A(N788), .B(N797), .CI(N790));
ADDFX1 inst_cellmath__62_0_I292 (.CO(inst_cellmath__62_0_out1[20]), .S(inst_cellmath__62_0_out0[19]), .A(N792), .B(N799), .CI(N801));
ADDFX1 inst_cellmath__62_0_I293 (.CO(N806), .S(N805), .A(N506), .B(N638), .CI(N572));
ADDFX1 inst_cellmath__62_0_I294 (.CO(N808), .S(N807), .A(N539), .B(N605), .CI(N796));
ADDFX1 inst_cellmath__62_0_I295 (.CO(N810), .S(N809), .A(N805), .B(N798), .CI(N807));
ADDFX1 inst_cellmath__62_0_I296 (.CO(inst_cellmath__62_0_out1[21]), .S(inst_cellmath__62_0_out0[20]), .A(N802), .B(N800), .CI(N809));
ADDFX1 inst_cellmath__62_0_I297 (.CO(N814), .S(N813), .A(N607), .B(N541), .CI(N640));
ADDFX1 inst_cellmath__62_0_I298 (.CO(N816), .S(N815), .A(N806), .B(N574), .CI(N813));
ADDFX1 inst_cellmath__62_0_I299 (.CO(inst_cellmath__62_0_out0[22]), .S(inst_cellmath__62_0_out0[21]), .A(N815), .B(N808), .CI(N810));
ADDFX1 inst_cellmath__62_0_I300 (.CO(N820), .S(N819), .A(N642), .B(N576), .CI(N609));
ADDFX1 inst_cellmath__62_0_I301 (.CO(inst_cellmath__62_0_out0[23]), .S(inst_cellmath__62_0_out1[22]), .A(N819), .B(N814), .CI(N816));
ADDFX1 inst_cellmath__62_0_I302 (.CO(inst_cellmath__62_0_out0[24]), .S(inst_cellmath__62_0_out1[23]), .A(N644), .B(N611), .CI(N820));
assign inst_cellmath__62_0_out0[0] = 1'B0;
assign inst_cellmath__62_0_out0[1] = 1'B0;
assign inst_cellmath__62_0_out0[2] = 1'B0;
assign inst_cellmath__62_0_out0[3] = 1'B0;
assign inst_cellmath__62_0_out0[4] = 1'B0;
assign inst_cellmath__62_0_out0[25] = 1'B0;
assign inst_cellmath__62_0_out0[26] = 1'B0;
assign inst_cellmath__62_0_out0[27] = 1'B0;
assign inst_cellmath__62_0_out0[28] = 1'B0;
assign inst_cellmath__62_0_out0[29] = 1'B0;
assign inst_cellmath__62_0_out0[30] = 1'B0;
assign inst_cellmath__62_0_out0[31] = 1'B0;
assign inst_cellmath__62_0_out0[32] = 1'B0;
assign inst_cellmath__62_0_out0[33] = 1'B0;
assign inst_cellmath__62_0_out0[34] = 1'B0;
assign inst_cellmath__62_0_out0[35] = 1'B0;
assign inst_cellmath__62_0_out0[36] = 1'B0;
assign inst_cellmath__62_0_out0[37] = 1'B0;
assign inst_cellmath__62_0_out0[38] = 1'B0;
assign inst_cellmath__62_0_out0[39] = 1'B0;
assign inst_cellmath__62_0_out1[0] = 1'B0;
assign inst_cellmath__62_0_out1[1] = 1'B0;
assign inst_cellmath__62_0_out1[2] = 1'B0;
assign inst_cellmath__62_0_out1[3] = 1'B0;
assign inst_cellmath__62_0_out1[25] = 1'B0;
assign inst_cellmath__62_0_out1[26] = 1'B0;
assign inst_cellmath__62_0_out1[27] = 1'B0;
assign inst_cellmath__62_0_out1[28] = 1'B0;
assign inst_cellmath__62_0_out1[29] = 1'B0;
assign inst_cellmath__62_0_out1[30] = 1'B0;
assign inst_cellmath__62_0_out1[31] = 1'B0;
assign inst_cellmath__62_0_out1[32] = 1'B0;
assign inst_cellmath__62_0_out1[33] = 1'B0;
assign inst_cellmath__62_0_out1[34] = 1'B0;
assign inst_cellmath__62_0_out1[35] = 1'B0;
assign inst_cellmath__62_0_out1[36] = 1'B0;
assign inst_cellmath__62_0_out1[37] = 1'B0;
assign inst_cellmath__62_0_out1[38] = 1'B0;
assign inst_cellmath__62_0_out1[39] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_cellmath__63_0_bdw1471647203_bdw (
	inst_cellmath__63_0_out0,
	inst_cellmath__63_0_out1,
	inst_cellmath__63_0_in0,
	inst_cellmath__63_0_in1,
	inst_cellmath__63_0_in2
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__63_0_out0,
	inst_cellmath__63_0_out1;
input [27:10] inst_cellmath__63_0_in0;
input  inst_cellmath__63_0_in1;
input [14:0] inst_cellmath__63_0_in2;
wire N414,N416,N418,N420,N422,N424,N426 
	,N428,N430,N432,N434,N436,N438,N440,N442 
	,N444,N462,N464,N466,N468,N470,N472,N474 
	,N476,N478,N480,N482,N484,N486,N488,N490 
	,N492,N506,N508,N510,N512,N514,N516,N518 
	,N520,N522,N524,N526,N528,N530,N532,N534 
	,N536,N538,N540,N554,N556,N558,N560,N562 
	,N564,N566,N568,N570,N572,N574,N576,N578 
	,N580,N582,N584,N586,N588,N602,N604,N606 
	,N608,N610,N612,N614,N616,N618,N620,N622 
	,N624,N626,N628,N630,N632,N634,N636,N650 
	,N652,N654,N656,N658,N660,N662,N664,N666 
	,N668,N670,N672,N674,N676,N678,N680,N682 
	,N684,N698,N700,N702,N704,N706,N708,N710 
	,N712,N714,N716,N718,N720,N722,N724,N726 
	,N728,N730,N732,N746,N748,N750,N752,N754 
	,N756,N758,N760,N762,N764,N766,N768,N770 
	,N772,N774,N776,N778,N780,N794,N796,N798 
	,N800,N802,N804,N806,N808,N810,N812,N814 
	,N816,N818,N820,N822,N824,N826,N828,N842 
	,N844,N846,N848,N850,N852,N854,N856,N858 
	,N860,N862,N864,N866,N868,N870,N872,N874 
	,N876,N890,N892,N894,N896,N898,N900,N902 
	,N904,N906,N908,N910,N912,N914,N916,N918 
	,N920,N922,N924,N938,N940,N942,N944,N946 
	,N948,N950,N952,N954,N956,N958,N960,N962 
	,N964,N966,N968,N970,N972,N986,N988,N990 
	,N992,N994,N996,N998,N1000,N1002,N1004,N1006 
	,N1008,N1010,N1012,N1014,N1016,N1018,N1020,N1034 
	,N1036,N1038,N1040,N1042,N1044,N1046,N1048,N1050 
	,N1052,N1054,N1056,N1058,N1060,N1062,N1064,N1066 
	,N1068,N1082,N1084,N1086,N1088,N1090,N1092,N1094 
	,N1096,N1098,N1100,N1102,N1104,N1106,N1108,N1110 
	,N1112,N1114,N1116,N1130,N1132,N1134,N1136,N1138 
	,N1140,N1142,N1144,N1146,N1148,N1150,N1152,N1154 
	,N1156,N1158,N1160,N1162,N1164,N1186,N1187,N1189 
	,N1190,N1191,N1193,N1196,N1197,N1198,N1199,N1200 
	,N1201,N1204,N1205,N1206,N1207,N1208,N1209,N1210 
	,N1211,N1214,N1215,N1216,N1217,N1218,N1219,N1220 
	,N1221,N1222,N1223,N1226,N1227,N1228,N1229,N1230 
	,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1240 
	,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248 
	,N1249,N1250,N1251,N1252,N1253,N1256,N1257,N1258 
	,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266 
	,N1267,N1268,N1269,N1270,N1271,N1274,N1275,N1276 
	,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284 
	,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1294 
	,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302 
	,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310 
	,N1311,N1312,N1313,N1316,N1317,N1318,N1319,N1320 
	,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328 
	,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336 
	,N1337,N1340,N1341,N1342,N1343,N1344,N1345,N1346 
	,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354 
	,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362 
	,N1363,N1366,N1367,N1370,N1371,N1372,N1373,N1374 
	,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382 
	,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390 
	,N1391,N1392,N1393,N1396,N1397,N1398,N1399,N1400 
	,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408 
	,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416 
	,N1417,N1418,N1419,N1420,N1421,N1424,N1425,N1426 
	,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434 
	,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442 
	,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1452 
	,N1453,N1456,N1457,N1458,N1459,N1460,N1461,N1462 
	,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470 
	,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478 
	,N1479,N1482,N1483,N1484,N1485,N1486,N1487,N1488 
	,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496 
	,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504 
	,N1505,N1506,N1507,N1510,N1511,N1512,N1513,N1514 
	,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522 
	,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530 
	,N1531,N1532,N1533,N1536,N1537,N1538,N1539,N1540 
	,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548 
	,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556 
	,N1557,N1560,N1561,N1562,N1563,N1564,N1565,N1566 
	,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574 
	,N1575,N1576,N1577,N1578,N1579,N1582,N1583,N1584 
	,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592 
	,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1602 
	,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610 
	,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1620 
	,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628 
	,N1629,N1630,N1631,N1632,N1633,N1636,N1637,N1638 
	,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646 
	,N1647,N1650,N1651,N1652,N1653,N1654,N1655,N1656 
	,N1657,N1658,N1659,N1662,N1663,N1664,N1665,N1666 
	,N1667,N1668,N1669,N1672,N1673,N1674,N1675,N1676 
	,N1677,N1680,N1681,N1682,N1683,N1686,N1687,N1803 
	,N1808,N1809,N1813,N1816,N1817,N1818,N1819,N1820 
	,N1821,N1822,N1823,N1825,N1826,N1827,N1828,N1829 
	,N1831,N1832,N1834,N1835,N1836,N1837,N1838,N1840 
	,N1841,N1843,N1844,N1847,N1849,N1850,N1852,N1853 
	,N1855,N1856,N1858,N1864,N1867,N1870,N1871,N1878 
	,N1885,N1892,N1899,N1906,N1913,N1920,N1921,N1922 
	,N1929,N1930,N1931,N1938,N1939;
BUFX3 inst_cellmath__63_0_I866 (.Y(N1808), .A(inst_cellmath__63_0_in0[10]));
CLKINVX4 inst_cellmath__63_0_I722 (.Y(N1809), .A(N1808));
BUFX2 inst_cellmath__63_0_I867 (.Y(N1813), .A(inst_cellmath__63_0_in0[11]));
INVX2 inst_cellmath__63_0_I730 (.Y(N1817), .A(N1813));
INVX2 inst_cellmath__63_0_I729 (.Y(N1816), .A(N1813));
INVX3 inst_cellmath__63_0_I731 (.Y(N1818), .A(inst_cellmath__63_0_in0[12]));
INVX3 inst_cellmath__63_0_I732 (.Y(N1819), .A(N1818));
CLKINVX4 inst_cellmath__63_0_I733 (.Y(N1820), .A(N1819));
INVX2 inst_cellmath__63_0_I734 (.Y(N1821), .A(inst_cellmath__63_0_in0[13]));
INVX3 inst_cellmath__63_0_I735 (.Y(N1822), .A(N1821));
INVX3 inst_cellmath__63_0_I736 (.Y(N1823), .A(N1822));
BUFX3 inst_cellmath__63_0_I870 (.Y(N1825), .A(inst_cellmath__63_0_in0[14]));
INVX3 inst_cellmath__63_0_I739 (.Y(N1826), .A(N1825));
INVX2 inst_cellmath__63_0_I740 (.Y(N1827), .A(inst_cellmath__63_0_in0[15]));
INVX3 inst_cellmath__63_0_I741 (.Y(N1828), .A(N1827));
INVX3 inst_cellmath__63_0_I742 (.Y(N1829), .A(N1828));
BUFX3 inst_cellmath__63_0_I872 (.Y(N1831), .A(inst_cellmath__63_0_in0[16]));
INVX3 inst_cellmath__63_0_I745 (.Y(N1832), .A(N1831));
BUFX3 inst_cellmath__63_0_I873 (.Y(N1834), .A(inst_cellmath__63_0_in0[17]));
INVX3 inst_cellmath__63_0_I748 (.Y(N1835), .A(N1834));
INVX2 inst_cellmath__63_0_I749 (.Y(N1836), .A(inst_cellmath__63_0_in0[18]));
INVX2 inst_cellmath__63_0_I750 (.Y(N1837), .A(N1836));
INVX3 inst_cellmath__63_0_I751 (.Y(N1838), .A(N1837));
BUFX3 inst_cellmath__63_0_I875 (.Y(N1840), .A(inst_cellmath__63_0_in0[19]));
INVX3 inst_cellmath__63_0_I754 (.Y(N1841), .A(N1840));
BUFX2 inst_cellmath__63_0_I876 (.Y(N1843), .A(inst_cellmath__63_0_in0[20]));
INVX3 inst_cellmath__63_0_I757 (.Y(N1844), .A(N1843));
INVX1 inst_cellmath__63_0_I760 (.Y(N1847), .A(inst_cellmath__63_0_in0[21]));
CLKBUFX12 inst_cellmath__63_0_I878 (.Y(N1849), .A(inst_cellmath__63_0_in0[22]));
INVX20 inst_cellmath__63_0_I763 (.Y(N1850), .A(N1849));
BUFX2 inst_cellmath__63_0_I879 (.Y(N1852), .A(inst_cellmath__63_0_in0[23]));
INVX3 inst_cellmath__63_0_I766 (.Y(N1853), .A(N1852));
BUFX3 inst_cellmath__63_0_I880 (.Y(N1855), .A(inst_cellmath__63_0_in0[24]));
CLKINVX4 inst_cellmath__63_0_I769 (.Y(N1856), .A(N1855));
CLKBUFX12 inst_cellmath__63_0_I881 (.Y(N1858), .A(inst_cellmath__63_0_in0[25]));
INVX20 inst_cellmath__63_0_I777 (.Y(N1864), .A(N1858));
INVX1 inst_cellmath__63_0_I780 (.Y(N1867), .A(inst_cellmath__63_0_in0[26]));
INVX1 inst_cellmath__63_0_I783 (.Y(N1870), .A(inst_cellmath__63_0_in0[27]));
INVXL inst_cellmath__63_0_I784 (.Y(N1871), .A(inst_cellmath__63_0_in2[0]));
NOR2XL inst_cellmath__63_0_I66 (.Y(inst_cellmath__63_0_out1[0]), .A(N1871), .B(N1809));
NOR2XL inst_cellmath__63_0_I67 (.Y(inst_cellmath__63_0_out0[1]), .A(N1871), .B(N1817));
NOR2XL inst_cellmath__63_0_I68 (.Y(N414), .A(N1871), .B(N1820));
NOR2X1 inst_cellmath__63_0_I69 (.Y(N416), .A(N1871), .B(N1823));
NOR2XL inst_cellmath__63_0_I70 (.Y(N418), .A(N1871), .B(N1826));
NOR2XL inst_cellmath__63_0_I71 (.Y(N420), .A(N1871), .B(N1829));
NOR2X1 inst_cellmath__63_0_I72 (.Y(N422), .A(N1871), .B(N1832));
NOR2XL inst_cellmath__63_0_I73 (.Y(N424), .A(N1871), .B(N1835));
NOR2XL inst_cellmath__63_0_I74 (.Y(N426), .A(N1871), .B(N1838));
NOR2XL inst_cellmath__63_0_I75 (.Y(N428), .A(N1871), .B(N1841));
NOR2XL inst_cellmath__63_0_I76 (.Y(N430), .A(N1871), .B(N1844));
NOR2XL inst_cellmath__63_0_I77 (.Y(N432), .A(N1871), .B(N1847));
NOR2X2 inst_cellmath__63_0_I78 (.Y(N434), .A(N1871), .B(N1850));
NOR2XL inst_cellmath__63_0_I79 (.Y(N436), .A(N1871), .B(N1853));
NOR2XL inst_cellmath__63_0_I80 (.Y(N438), .A(N1871), .B(N1856));
NOR2X2 inst_cellmath__63_0_I81 (.Y(N440), .A(N1871), .B(N1864));
NOR2XL inst_cellmath__63_0_I82 (.Y(N442), .A(N1871), .B(N1867));
NOR2XL inst_cellmath__63_0_I83 (.Y(N444), .A(N1871), .B(N1870));
INVXL inst_cellmath__63_0_I791 (.Y(N1878), .A(inst_cellmath__63_0_in2[1]));
NOR2XL inst_cellmath__63_0_I89 (.Y(inst_cellmath__63_0_out1[1]), .A(N1878), .B(N1809));
NOR2XL inst_cellmath__63_0_I90 (.Y(inst_cellmath__63_0_out1[2]), .A(N1878), .B(N1817));
NOR2X2 inst_cellmath__63_0_I91 (.Y(N462), .A(N1878), .B(N1820));
NOR2XL inst_cellmath__63_0_I92 (.Y(N464), .A(N1878), .B(N1823));
NOR2XL inst_cellmath__63_0_I93 (.Y(N466), .A(N1878), .B(N1826));
NOR2XL inst_cellmath__63_0_I94 (.Y(N468), .A(N1878), .B(N1829));
NOR2XL inst_cellmath__63_0_I95 (.Y(N470), .A(N1878), .B(N1832));
NOR2XL inst_cellmath__63_0_I96 (.Y(N472), .A(N1878), .B(N1835));
NOR2XL inst_cellmath__63_0_I97 (.Y(N474), .A(N1878), .B(N1838));
NOR2XL inst_cellmath__63_0_I98 (.Y(N476), .A(N1878), .B(N1841));
NOR2XL inst_cellmath__63_0_I99 (.Y(N478), .A(N1878), .B(N1844));
NOR2XL inst_cellmath__63_0_I100 (.Y(N480), .A(N1878), .B(N1847));
NOR2XL inst_cellmath__63_0_I101 (.Y(N482), .A(N1878), .B(N1850));
NOR2XL inst_cellmath__63_0_I102 (.Y(N484), .A(N1878), .B(N1853));
NOR2XL inst_cellmath__63_0_I103 (.Y(N486), .A(N1878), .B(N1856));
NOR2X2 inst_cellmath__63_0_I104 (.Y(N488), .A(N1878), .B(N1864));
NOR2XL inst_cellmath__63_0_I105 (.Y(N490), .A(N1878), .B(N1867));
NOR2XL inst_cellmath__63_0_I106 (.Y(N492), .A(N1878), .B(N1870));
INVXL inst_cellmath__63_0_I798 (.Y(N1885), .A(inst_cellmath__63_0_in2[2]));
NOR2XL inst_cellmath__63_0_I112 (.Y(N506), .A(N1885), .B(N1809));
NOR2X1 inst_cellmath__63_0_I113 (.Y(N508), .A(N1885), .B(N1817));
NOR2XL inst_cellmath__63_0_I114 (.Y(N510), .A(N1885), .B(N1820));
NOR2XL inst_cellmath__63_0_I115 (.Y(N512), .A(N1885), .B(N1823));
NOR2XL inst_cellmath__63_0_I116 (.Y(N514), .A(N1885), .B(N1826));
NOR2XL inst_cellmath__63_0_I117 (.Y(N516), .A(N1885), .B(N1829));
NOR2XL inst_cellmath__63_0_I118 (.Y(N518), .A(N1885), .B(N1832));
NOR2XL inst_cellmath__63_0_I119 (.Y(N520), .A(N1885), .B(N1835));
NOR2XL inst_cellmath__63_0_I120 (.Y(N522), .A(N1885), .B(N1838));
NOR2XL inst_cellmath__63_0_I121 (.Y(N524), .A(N1885), .B(N1841));
NOR2XL inst_cellmath__63_0_I122 (.Y(N526), .A(N1885), .B(N1844));
NOR2XL inst_cellmath__63_0_I123 (.Y(N528), .A(N1885), .B(N1847));
NOR2XL inst_cellmath__63_0_I124 (.Y(N530), .A(N1885), .B(N1850));
NOR2X1 inst_cellmath__63_0_I125 (.Y(N532), .A(N1885), .B(N1853));
NOR2XL inst_cellmath__63_0_I126 (.Y(N534), .A(N1885), .B(N1856));
NOR2X2 inst_cellmath__63_0_I127 (.Y(N536), .A(N1885), .B(N1864));
NOR2XL inst_cellmath__63_0_I128 (.Y(N538), .A(N1885), .B(N1867));
NOR2XL inst_cellmath__63_0_I129 (.Y(N540), .A(N1885), .B(N1870));
INVXL inst_cellmath__63_0_I805 (.Y(N1892), .A(inst_cellmath__63_0_in2[3]));
NOR2X1 inst_cellmath__63_0_I135 (.Y(N554), .A(N1892), .B(N1809));
NOR2XL inst_cellmath__63_0_I136 (.Y(N556), .A(N1892), .B(N1816));
NOR2XL inst_cellmath__63_0_I137 (.Y(N558), .A(N1892), .B(N1820));
NOR2X2 inst_cellmath__63_0_I138 (.Y(N560), .A(N1892), .B(N1823));
NOR2X1 inst_cellmath__63_0_I139 (.Y(N562), .A(N1892), .B(N1826));
NOR2XL inst_cellmath__63_0_I140 (.Y(N564), .A(N1892), .B(N1829));
NOR2XL inst_cellmath__63_0_I141 (.Y(N566), .A(N1892), .B(N1832));
NOR2XL inst_cellmath__63_0_I142 (.Y(N568), .A(N1892), .B(N1835));
NOR2XL inst_cellmath__63_0_I143 (.Y(N570), .A(N1892), .B(N1838));
NOR2XL inst_cellmath__63_0_I144 (.Y(N572), .A(N1892), .B(N1841));
NOR2XL inst_cellmath__63_0_I145 (.Y(N574), .A(N1892), .B(N1844));
NOR2XL inst_cellmath__63_0_I146 (.Y(N576), .A(N1892), .B(N1847));
NOR2XL inst_cellmath__63_0_I147 (.Y(N578), .A(N1892), .B(N1850));
NOR2X1 inst_cellmath__63_0_I148 (.Y(N580), .A(N1892), .B(N1853));
NOR2XL inst_cellmath__63_0_I149 (.Y(N582), .A(N1892), .B(N1856));
NOR2X1 inst_cellmath__63_0_I150 (.Y(N584), .A(N1892), .B(N1864));
NOR2XL inst_cellmath__63_0_I151 (.Y(N586), .A(N1892), .B(N1867));
NOR2XL inst_cellmath__63_0_I152 (.Y(N588), .A(N1892), .B(N1870));
INVXL inst_cellmath__63_0_I812 (.Y(N1899), .A(inst_cellmath__63_0_in2[4]));
NOR2XL inst_cellmath__63_0_I158 (.Y(N602), .A(N1899), .B(N1809));
NOR2XL inst_cellmath__63_0_I159 (.Y(N604), .A(N1899), .B(N1816));
NOR2X1 inst_cellmath__63_0_I160 (.Y(N606), .A(N1899), .B(N1820));
NOR2XL inst_cellmath__63_0_I161 (.Y(N608), .A(N1899), .B(N1823));
NOR2X1 inst_cellmath__63_0_I162 (.Y(N610), .A(N1899), .B(N1826));
NOR2XL inst_cellmath__63_0_I163 (.Y(N612), .A(N1899), .B(N1829));
NOR2XL inst_cellmath__63_0_I164 (.Y(N614), .A(N1899), .B(N1832));
NOR2XL inst_cellmath__63_0_I165 (.Y(N616), .A(N1899), .B(N1835));
NOR2XL inst_cellmath__63_0_I166 (.Y(N618), .A(N1899), .B(N1838));
NOR2XL inst_cellmath__63_0_I167 (.Y(N620), .A(N1899), .B(N1841));
NOR2XL inst_cellmath__63_0_I168 (.Y(N622), .A(N1899), .B(N1844));
NOR2XL inst_cellmath__63_0_I169 (.Y(N624), .A(N1899), .B(N1847));
NOR2XL inst_cellmath__63_0_I170 (.Y(N626), .A(N1899), .B(N1850));
NOR2XL inst_cellmath__63_0_I171 (.Y(N628), .A(N1899), .B(N1853));
NOR2XL inst_cellmath__63_0_I172 (.Y(N630), .A(N1899), .B(N1856));
NOR2X1 inst_cellmath__63_0_I173 (.Y(N632), .A(N1899), .B(N1864));
NOR2XL inst_cellmath__63_0_I174 (.Y(N634), .A(N1899), .B(N1867));
NOR2XL inst_cellmath__63_0_I175 (.Y(N636), .A(N1899), .B(N1870));
INVXL inst_cellmath__63_0_I819 (.Y(N1906), .A(inst_cellmath__63_0_in2[5]));
NOR2X1 inst_cellmath__63_0_I181 (.Y(N650), .A(N1906), .B(N1809));
NOR2XL inst_cellmath__63_0_I182 (.Y(N652), .A(N1906), .B(N1816));
NOR2XL inst_cellmath__63_0_I183 (.Y(N654), .A(N1906), .B(N1820));
NOR2XL inst_cellmath__63_0_I184 (.Y(N656), .A(N1906), .B(N1823));
NOR2XL inst_cellmath__63_0_I185 (.Y(N658), .A(N1906), .B(N1826));
NOR2XL inst_cellmath__63_0_I186 (.Y(N660), .A(N1906), .B(N1829));
NOR2XL inst_cellmath__63_0_I187 (.Y(N662), .A(N1906), .B(N1832));
NOR2XL inst_cellmath__63_0_I188 (.Y(N664), .A(N1906), .B(N1835));
NOR2XL inst_cellmath__63_0_I189 (.Y(N666), .A(N1906), .B(N1838));
NOR2XL inst_cellmath__63_0_I190 (.Y(N668), .A(N1906), .B(N1841));
NOR2XL inst_cellmath__63_0_I191 (.Y(N670), .A(N1906), .B(N1844));
NOR2XL inst_cellmath__63_0_I192 (.Y(N672), .A(N1906), .B(N1847));
NOR2XL inst_cellmath__63_0_I193 (.Y(N674), .A(N1906), .B(N1850));
NOR2XL inst_cellmath__63_0_I194 (.Y(N676), .A(N1906), .B(N1853));
NOR2XL inst_cellmath__63_0_I195 (.Y(N678), .A(N1906), .B(N1856));
NOR2XL inst_cellmath__63_0_I196 (.Y(N680), .A(N1906), .B(N1864));
NOR2XL inst_cellmath__63_0_I197 (.Y(N682), .A(N1906), .B(N1867));
NOR2XL inst_cellmath__63_0_I198 (.Y(N684), .A(N1906), .B(N1870));
INVXL inst_cellmath__63_0_I826 (.Y(N1913), .A(inst_cellmath__63_0_in2[6]));
NOR2XL inst_cellmath__63_0_I204 (.Y(N698), .A(N1913), .B(N1809));
NOR2XL inst_cellmath__63_0_I205 (.Y(N700), .A(N1913), .B(N1816));
NOR2XL inst_cellmath__63_0_I206 (.Y(N702), .A(N1913), .B(N1820));
NOR2XL inst_cellmath__63_0_I207 (.Y(N704), .A(N1913), .B(N1823));
NOR2XL inst_cellmath__63_0_I208 (.Y(N706), .A(N1913), .B(N1826));
NOR2XL inst_cellmath__63_0_I209 (.Y(N708), .A(N1913), .B(N1829));
NOR2XL inst_cellmath__63_0_I210 (.Y(N710), .A(N1913), .B(N1832));
NOR2XL inst_cellmath__63_0_I211 (.Y(N712), .A(N1913), .B(N1835));
NOR2XL inst_cellmath__63_0_I212 (.Y(N714), .A(N1913), .B(N1838));
NOR2XL inst_cellmath__63_0_I213 (.Y(N716), .A(N1913), .B(N1841));
NOR2XL inst_cellmath__63_0_I214 (.Y(N718), .A(N1913), .B(N1844));
NOR2XL inst_cellmath__63_0_I215 (.Y(N720), .A(N1913), .B(N1847));
NOR2XL inst_cellmath__63_0_I216 (.Y(N722), .A(N1913), .B(N1850));
NOR2XL inst_cellmath__63_0_I217 (.Y(N724), .A(N1913), .B(N1853));
NOR2XL inst_cellmath__63_0_I218 (.Y(N726), .A(N1913), .B(N1856));
NOR2XL inst_cellmath__63_0_I219 (.Y(N728), .A(N1913), .B(N1864));
NOR2XL inst_cellmath__63_0_I220 (.Y(N730), .A(N1913), .B(N1867));
NOR2XL inst_cellmath__63_0_I221 (.Y(N732), .A(N1913), .B(N1870));
INVXL inst_cellmath__63_0_I833 (.Y(N1920), .A(inst_cellmath__63_0_in2[7]));
NOR2X1 inst_cellmath__63_0_I227 (.Y(N746), .A(N1920), .B(N1809));
NOR2XL inst_cellmath__63_0_I228 (.Y(N748), .A(N1920), .B(N1816));
NOR2XL inst_cellmath__63_0_I229 (.Y(N750), .A(N1920), .B(N1820));
NOR2X1 inst_cellmath__63_0_I230 (.Y(N752), .A(N1920), .B(N1823));
NOR2XL inst_cellmath__63_0_I231 (.Y(N754), .A(N1920), .B(N1826));
NOR2XL inst_cellmath__63_0_I232 (.Y(N756), .A(N1920), .B(N1829));
NOR2XL inst_cellmath__63_0_I233 (.Y(N758), .A(N1920), .B(N1832));
NOR2XL inst_cellmath__63_0_I234 (.Y(N760), .A(N1920), .B(N1835));
NOR2XL inst_cellmath__63_0_I235 (.Y(N762), .A(N1920), .B(N1838));
NOR2XL inst_cellmath__63_0_I236 (.Y(N764), .A(N1920), .B(N1841));
NOR2XL inst_cellmath__63_0_I237 (.Y(N766), .A(N1920), .B(N1844));
NOR2XL inst_cellmath__63_0_I238 (.Y(N768), .A(N1920), .B(N1847));
NOR2XL inst_cellmath__63_0_I239 (.Y(N770), .A(N1920), .B(N1850));
NOR2XL inst_cellmath__63_0_I240 (.Y(N772), .A(N1920), .B(N1853));
NOR2XL inst_cellmath__63_0_I241 (.Y(N774), .A(N1920), .B(N1856));
NOR2XL inst_cellmath__63_0_I242 (.Y(N776), .A(N1920), .B(N1864));
NOR2XL inst_cellmath__63_0_I243 (.Y(N778), .A(N1920), .B(N1867));
NOR2XL inst_cellmath__63_0_I244 (.Y(N780), .A(N1920), .B(N1870));
INVXL inst_cellmath__63_0_I834 (.Y(N1921), .A(inst_cellmath__63_0_in2[8]));
NOR2XL inst_cellmath__63_0_I250 (.Y(N794), .A(N1921), .B(N1809));
NOR2XL inst_cellmath__63_0_I251 (.Y(N796), .A(N1921), .B(N1816));
NOR2XL inst_cellmath__63_0_I252 (.Y(N798), .A(N1921), .B(N1820));
NOR2XL inst_cellmath__63_0_I253 (.Y(N800), .A(N1921), .B(N1823));
NOR2XL inst_cellmath__63_0_I254 (.Y(N802), .A(N1921), .B(N1826));
NOR2XL inst_cellmath__63_0_I255 (.Y(N804), .A(N1921), .B(N1829));
NOR2XL inst_cellmath__63_0_I256 (.Y(N806), .A(N1921), .B(N1832));
NOR2XL inst_cellmath__63_0_I257 (.Y(N808), .A(N1921), .B(N1835));
NOR2XL inst_cellmath__63_0_I258 (.Y(N810), .A(N1921), .B(N1838));
NOR2XL inst_cellmath__63_0_I259 (.Y(N812), .A(N1921), .B(N1841));
NOR2XL inst_cellmath__63_0_I260 (.Y(N814), .A(N1921), .B(N1844));
NOR2XL inst_cellmath__63_0_I261 (.Y(N816), .A(N1921), .B(N1847));
NOR2XL inst_cellmath__63_0_I262 (.Y(N818), .A(N1921), .B(N1850));
NOR2XL inst_cellmath__63_0_I263 (.Y(N820), .A(N1921), .B(N1853));
NOR2XL inst_cellmath__63_0_I264 (.Y(N822), .A(N1921), .B(N1856));
NOR2XL inst_cellmath__63_0_I265 (.Y(N824), .A(N1921), .B(N1864));
NOR2XL inst_cellmath__63_0_I266 (.Y(N826), .A(N1921), .B(N1867));
NOR2XL inst_cellmath__63_0_I267 (.Y(N828), .A(N1921), .B(N1870));
INVXL inst_cellmath__63_0_I835 (.Y(N1922), .A(inst_cellmath__63_0_in2[9]));
NOR2XL inst_cellmath__63_0_I273 (.Y(N842), .A(N1922), .B(N1809));
NOR2XL inst_cellmath__63_0_I274 (.Y(N844), .A(N1922), .B(N1816));
NOR2XL inst_cellmath__63_0_I275 (.Y(N846), .A(N1922), .B(N1820));
NOR2XL inst_cellmath__63_0_I276 (.Y(N848), .A(N1922), .B(N1823));
NOR2XL inst_cellmath__63_0_I277 (.Y(N850), .A(N1922), .B(N1826));
NOR2XL inst_cellmath__63_0_I278 (.Y(N852), .A(N1922), .B(N1829));
NOR2XL inst_cellmath__63_0_I279 (.Y(N854), .A(N1922), .B(N1832));
NOR2XL inst_cellmath__63_0_I280 (.Y(N856), .A(N1922), .B(N1835));
NOR2XL inst_cellmath__63_0_I281 (.Y(N858), .A(N1922), .B(N1838));
NOR2X1 inst_cellmath__63_0_I282 (.Y(N860), .A(N1922), .B(N1841));
NOR2XL inst_cellmath__63_0_I283 (.Y(N862), .A(N1922), .B(N1844));
NOR2XL inst_cellmath__63_0_I284 (.Y(N864), .A(N1922), .B(N1847));
NOR2XL inst_cellmath__63_0_I285 (.Y(N866), .A(N1922), .B(N1850));
NOR2XL inst_cellmath__63_0_I286 (.Y(N868), .A(N1922), .B(N1853));
NOR2XL inst_cellmath__63_0_I287 (.Y(N870), .A(N1922), .B(N1856));
NOR2XL inst_cellmath__63_0_I288 (.Y(N872), .A(N1922), .B(N1864));
NOR2XL inst_cellmath__63_0_I289 (.Y(N874), .A(N1922), .B(N1867));
NOR2XL inst_cellmath__63_0_I290 (.Y(N876), .A(N1922), .B(N1870));
INVXL inst_cellmath__63_0_I842 (.Y(N1929), .A(inst_cellmath__63_0_in2[10]));
NOR2XL inst_cellmath__63_0_I296 (.Y(N890), .A(N1929), .B(N1809));
NOR2XL inst_cellmath__63_0_I297 (.Y(N892), .A(N1929), .B(N1816));
NOR2XL inst_cellmath__63_0_I298 (.Y(N894), .A(N1929), .B(N1820));
NOR2XL inst_cellmath__63_0_I299 (.Y(N896), .A(N1929), .B(N1823));
NOR2XL inst_cellmath__63_0_I300 (.Y(N898), .A(N1929), .B(N1826));
NOR2XL inst_cellmath__63_0_I301 (.Y(N900), .A(N1929), .B(N1829));
NOR2XL inst_cellmath__63_0_I302 (.Y(N902), .A(N1929), .B(N1832));
NOR2X1 inst_cellmath__63_0_I303 (.Y(N904), .A(N1929), .B(N1835));
NOR2XL inst_cellmath__63_0_I304 (.Y(N906), .A(N1929), .B(N1838));
NOR2XL inst_cellmath__63_0_I305 (.Y(N908), .A(N1929), .B(N1841));
NOR2XL inst_cellmath__63_0_I306 (.Y(N910), .A(N1929), .B(N1844));
NOR2XL inst_cellmath__63_0_I307 (.Y(N912), .A(N1929), .B(N1847));
NOR2XL inst_cellmath__63_0_I308 (.Y(N914), .A(N1929), .B(N1850));
NOR2XL inst_cellmath__63_0_I309 (.Y(N916), .A(N1929), .B(N1853));
NOR2XL inst_cellmath__63_0_I310 (.Y(N918), .A(N1929), .B(N1856));
NOR2XL inst_cellmath__63_0_I311 (.Y(N920), .A(N1929), .B(N1864));
NOR2XL inst_cellmath__63_0_I312 (.Y(N922), .A(N1929), .B(N1867));
NOR2XL inst_cellmath__63_0_I313 (.Y(N924), .A(N1929), .B(N1870));
INVXL inst_cellmath__63_0_I843 (.Y(N1930), .A(inst_cellmath__63_0_in2[11]));
NOR2XL inst_cellmath__63_0_I319 (.Y(N938), .A(N1930), .B(N1809));
NOR2XL inst_cellmath__63_0_I320 (.Y(N940), .A(N1930), .B(N1817));
NOR2XL inst_cellmath__63_0_I321 (.Y(N942), .A(N1930), .B(N1820));
NOR2XL inst_cellmath__63_0_I322 (.Y(N944), .A(N1930), .B(N1823));
NOR2XL inst_cellmath__63_0_I323 (.Y(N946), .A(N1930), .B(N1826));
NOR2XL inst_cellmath__63_0_I324 (.Y(N948), .A(N1930), .B(N1829));
NOR2X1 inst_cellmath__63_0_I325 (.Y(N950), .A(N1930), .B(N1832));
NOR2XL inst_cellmath__63_0_I326 (.Y(N952), .A(N1930), .B(N1835));
NOR2XL inst_cellmath__63_0_I327 (.Y(N954), .A(N1930), .B(N1838));
NOR2XL inst_cellmath__63_0_I328 (.Y(N956), .A(N1930), .B(N1841));
NOR2XL inst_cellmath__63_0_I329 (.Y(N958), .A(N1930), .B(N1844));
NOR2XL inst_cellmath__63_0_I330 (.Y(N960), .A(N1930), .B(N1847));
NOR2XL inst_cellmath__63_0_I331 (.Y(N962), .A(N1930), .B(N1850));
NOR2XL inst_cellmath__63_0_I332 (.Y(N964), .A(N1930), .B(N1853));
NOR2XL inst_cellmath__63_0_I333 (.Y(N966), .A(N1930), .B(N1856));
NOR2XL inst_cellmath__63_0_I334 (.Y(N968), .A(N1930), .B(N1864));
NOR2XL inst_cellmath__63_0_I335 (.Y(N970), .A(N1930), .B(N1867));
NOR2XL inst_cellmath__63_0_I336 (.Y(N972), .A(N1930), .B(N1870));
INVXL inst_cellmath__63_0_I844 (.Y(N1931), .A(inst_cellmath__63_0_in2[12]));
NOR2XL inst_cellmath__63_0_I342 (.Y(N986), .A(N1931), .B(N1809));
NOR2XL inst_cellmath__63_0_I343 (.Y(N988), .A(N1931), .B(N1817));
NOR2XL inst_cellmath__63_0_I344 (.Y(N990), .A(N1931), .B(N1820));
NOR2XL inst_cellmath__63_0_I345 (.Y(N992), .A(N1931), .B(N1823));
NOR2X1 inst_cellmath__63_0_I346 (.Y(N994), .A(N1931), .B(N1826));
NOR2XL inst_cellmath__63_0_I347 (.Y(N996), .A(N1931), .B(N1829));
NOR2XL inst_cellmath__63_0_I348 (.Y(N998), .A(N1931), .B(N1832));
NOR2X1 inst_cellmath__63_0_I349 (.Y(N1000), .A(N1931), .B(N1835));
NOR2XL inst_cellmath__63_0_I350 (.Y(N1002), .A(N1931), .B(N1838));
NOR2XL inst_cellmath__63_0_I351 (.Y(N1004), .A(N1931), .B(N1841));
NOR2XL inst_cellmath__63_0_I352 (.Y(N1006), .A(N1931), .B(N1844));
NOR2XL inst_cellmath__63_0_I353 (.Y(N1008), .A(N1931), .B(N1847));
NOR2XL inst_cellmath__63_0_I354 (.Y(N1010), .A(N1931), .B(N1850));
NOR2XL inst_cellmath__63_0_I355 (.Y(N1012), .A(N1931), .B(N1853));
NOR2XL inst_cellmath__63_0_I356 (.Y(N1014), .A(N1931), .B(N1856));
NOR2XL inst_cellmath__63_0_I357 (.Y(N1016), .A(N1931), .B(N1864));
NOR2XL inst_cellmath__63_0_I358 (.Y(N1018), .A(N1931), .B(N1867));
NOR2XL inst_cellmath__63_0_I359 (.Y(N1020), .A(N1931), .B(N1870));
INVXL inst_cellmath__63_0_I851 (.Y(N1938), .A(inst_cellmath__63_0_in2[13]));
NOR2XL inst_cellmath__63_0_I365 (.Y(N1034), .A(N1938), .B(N1809));
NOR2XL inst_cellmath__63_0_I366 (.Y(N1036), .A(N1938), .B(N1817));
NOR2XL inst_cellmath__63_0_I367 (.Y(N1038), .A(N1938), .B(N1820));
NOR2XL inst_cellmath__63_0_I368 (.Y(N1040), .A(N1938), .B(N1823));
NOR2X1 inst_cellmath__63_0_I369 (.Y(N1042), .A(N1938), .B(N1826));
NOR2XL inst_cellmath__63_0_I370 (.Y(N1044), .A(N1938), .B(N1829));
NOR2XL inst_cellmath__63_0_I371 (.Y(N1046), .A(N1938), .B(N1832));
NOR2XL inst_cellmath__63_0_I372 (.Y(N1048), .A(N1938), .B(N1835));
NOR2XL inst_cellmath__63_0_I373 (.Y(N1050), .A(N1938), .B(N1838));
NOR2XL inst_cellmath__63_0_I374 (.Y(N1052), .A(N1938), .B(N1841));
NOR2XL inst_cellmath__63_0_I375 (.Y(N1054), .A(N1938), .B(N1844));
NOR2XL inst_cellmath__63_0_I376 (.Y(N1056), .A(N1938), .B(N1847));
NOR2XL inst_cellmath__63_0_I377 (.Y(N1058), .A(N1938), .B(N1850));
NOR2XL inst_cellmath__63_0_I378 (.Y(N1060), .A(N1938), .B(N1853));
NOR2XL inst_cellmath__63_0_I379 (.Y(N1062), .A(N1938), .B(N1856));
NOR2XL inst_cellmath__63_0_I380 (.Y(N1064), .A(N1938), .B(N1864));
NOR2XL inst_cellmath__63_0_I381 (.Y(N1066), .A(N1938), .B(N1867));
NOR2XL inst_cellmath__63_0_I382 (.Y(N1068), .A(N1938), .B(N1870));
INVXL inst_cellmath__63_0_I852 (.Y(N1939), .A(inst_cellmath__63_0_in2[14]));
NOR2X1 inst_cellmath__63_0_I388 (.Y(N1082), .A(N1939), .B(N1809));
NOR2XL inst_cellmath__63_0_I389 (.Y(N1084), .A(N1939), .B(N1817));
NOR2XL inst_cellmath__63_0_I390 (.Y(N1086), .A(N1939), .B(N1820));
NOR2XL inst_cellmath__63_0_I391 (.Y(N1088), .A(N1939), .B(N1823));
NOR2XL inst_cellmath__63_0_I392 (.Y(N1090), .A(N1939), .B(N1826));
NOR2X1 inst_cellmath__63_0_I393 (.Y(N1092), .A(N1939), .B(N1829));
NOR2XL inst_cellmath__63_0_I394 (.Y(N1094), .A(N1939), .B(N1832));
NOR2XL inst_cellmath__63_0_I395 (.Y(N1096), .A(N1939), .B(N1835));
NOR2XL inst_cellmath__63_0_I396 (.Y(N1098), .A(N1939), .B(N1838));
NOR2XL inst_cellmath__63_0_I397 (.Y(N1100), .A(N1939), .B(N1841));
NOR2XL inst_cellmath__63_0_I398 (.Y(N1102), .A(N1939), .B(N1844));
NOR2XL inst_cellmath__63_0_I399 (.Y(N1104), .A(N1939), .B(N1847));
NOR2XL inst_cellmath__63_0_I400 (.Y(N1106), .A(N1939), .B(N1850));
NOR2XL inst_cellmath__63_0_I401 (.Y(N1108), .A(N1939), .B(N1853));
NOR2XL inst_cellmath__63_0_I402 (.Y(N1110), .A(N1939), .B(N1856));
NOR2XL inst_cellmath__63_0_I403 (.Y(N1112), .A(N1939), .B(N1864));
NOR2XL inst_cellmath__63_0_I404 (.Y(N1114), .A(N1939), .B(N1867));
NOR2XL inst_cellmath__63_0_I405 (.Y(N1116), .A(N1939), .B(N1870));
BUFX3 inst_cellmath__63_0_I884 (.Y(inst_cellmath__63_0_out1[33]), .A(inst_cellmath__63_0_in1));
NAND2XL inst_cellmath__63_0_I411 (.Y(N1130), .A(inst_cellmath__63_0_out1[33]), .B(N1808));
NAND2X1 inst_cellmath__63_0_I412 (.Y(N1132), .A(inst_cellmath__63_0_out1[33]), .B(inst_cellmath__63_0_in0[11]));
NAND2XL inst_cellmath__63_0_I413 (.Y(N1134), .A(inst_cellmath__63_0_out1[33]), .B(N1819));
NAND2XL inst_cellmath__63_0_I414 (.Y(N1136), .A(inst_cellmath__63_0_out1[33]), .B(N1822));
NAND2X1 inst_cellmath__63_0_I415 (.Y(N1138), .A(inst_cellmath__63_0_out1[33]), .B(N1825));
NAND2X2 inst_cellmath__63_0_I416 (.Y(N1140), .A(inst_cellmath__63_0_out1[33]), .B(N1828));
NAND2XL inst_cellmath__63_0_I417 (.Y(N1142), .A(inst_cellmath__63_0_out1[33]), .B(N1831));
NAND2XL inst_cellmath__63_0_I418 (.Y(N1144), .A(inst_cellmath__63_0_out1[33]), .B(N1834));
NAND2XL inst_cellmath__63_0_I419 (.Y(N1146), .A(inst_cellmath__63_0_out1[33]), .B(N1837));
NAND2XL inst_cellmath__63_0_I420 (.Y(N1148), .A(inst_cellmath__63_0_out1[33]), .B(N1840));
NAND2XL inst_cellmath__63_0_I421 (.Y(N1150), .A(inst_cellmath__63_0_out1[33]), .B(N1843));
NAND2XL inst_cellmath__63_0_I422 (.Y(N1152), .A(inst_cellmath__63_0_out1[33]), .B(inst_cellmath__63_0_in0[21]));
NAND2XL inst_cellmath__63_0_I423 (.Y(N1154), .A(inst_cellmath__63_0_out1[33]), .B(N1849));
NAND2XL inst_cellmath__63_0_I424 (.Y(N1156), .A(inst_cellmath__63_0_out1[33]), .B(N1852));
NAND2XL inst_cellmath__63_0_I425 (.Y(N1158), .A(inst_cellmath__63_0_out1[33]), .B(N1855));
NAND2XL inst_cellmath__63_0_I426 (.Y(N1160), .A(inst_cellmath__63_0_out1[33]), .B(N1858));
NAND2XL inst_cellmath__63_0_I427 (.Y(N1162), .A(inst_cellmath__63_0_out1[33]), .B(inst_cellmath__63_0_in0[26]));
NAND2XL inst_cellmath__63_0_I428 (.Y(N1164), .A(inst_cellmath__63_0_out1[33]), .B(inst_cellmath__63_0_in0[27]));
ADDHX1 inst_cellmath__63_0_I446 (.CO(inst_cellmath__63_0_out1[3]), .S(inst_cellmath__63_0_out0[2]), .A(N414), .B(N506));
ADDHXL inst_cellmath__63_0_I447 (.CO(N1187), .S(N1186), .A(N462), .B(N416));
ADDFXL inst_cellmath__63_0_I448 (.CO(N1189), .S(inst_cellmath__63_0_out0[3]), .A(N508), .B(N554), .CI(N1186));
ADDHX1 inst_cellmath__63_0_I449 (.CO(N1191), .S(N1190), .A(N510), .B(N418));
ADDFX1 inst_cellmath__63_0_I450 (.CO(N1193), .S(inst_cellmath__63_0_out1[4]), .A(N602), .B(N464), .CI(N556));
ADDFXL inst_cellmath__63_0_I451 (.CO(inst_cellmath__63_0_out1[5]), .S(inst_cellmath__63_0_out0[4]), .A(N1190), .B(N1187), .CI(N1189));
ADDHX1 inst_cellmath__63_0_I452 (.CO(N1197), .S(N1196), .A(N420), .B(N466));
ADDFX1 inst_cellmath__63_0_I453 (.CO(N1199), .S(N1198), .A(N512), .B(N558), .CI(N650));
ADDFX1 inst_cellmath__63_0_I454 (.CO(N1201), .S(N1200), .A(N1191), .B(N604), .CI(N1196));
ADDFX1 inst_cellmath__63_0_I455 (.CO(inst_cellmath__63_0_out1[6]), .S(inst_cellmath__63_0_out0[5]), .A(N1198), .B(N1193), .CI(N1200));
ADDHX1 inst_cellmath__63_0_I456 (.CO(N1205), .S(N1204), .A(N468), .B(N514));
ADDFXL inst_cellmath__63_0_I457 (.CO(N1207), .S(N1206), .A(N560), .B(N606), .CI(N422));
ADDFX1 inst_cellmath__63_0_I458 (.CO(N1209), .S(N1208), .A(N652), .B(N698), .CI(N1197));
ADDFXL inst_cellmath__63_0_I459 (.CO(N1211), .S(N1210), .A(N1199), .B(N1204), .CI(N1206));
ADDFXL inst_cellmath__63_0_I460 (.CO(inst_cellmath__63_0_out1[7]), .S(inst_cellmath__63_0_out0[6]), .A(N1208), .B(N1201), .CI(N1210));
ADDHX1 inst_cellmath__63_0_I461 (.CO(N1215), .S(N1214), .A(N516), .B(N562));
ADDFX1 inst_cellmath__63_0_I462 (.CO(N1217), .S(N1216), .A(N608), .B(N654), .CI(N470));
ADDFX1 inst_cellmath__63_0_I463 (.CO(N1219), .S(N1218), .A(N746), .B(N424), .CI(N700));
ADDFX1 inst_cellmath__63_0_I464 (.CO(N1221), .S(N1220), .A(N1214), .B(N1205), .CI(N1207));
ADDFXL inst_cellmath__63_0_I465 (.CO(N1223), .S(N1222), .A(N1209), .B(N1216), .CI(N1218));
ADDFXL inst_cellmath__63_0_I466 (.CO(inst_cellmath__63_0_out1[8]), .S(inst_cellmath__63_0_out0[7]), .A(N1211), .B(N1220), .CI(N1222));
ADDHX1 inst_cellmath__63_0_I467 (.CO(N1227), .S(N1226), .A(N564), .B(N610));
ADDFX1 inst_cellmath__63_0_I468 (.CO(N1229), .S(N1228), .A(N656), .B(N702), .CI(N518));
ADDFX1 inst_cellmath__63_0_I469 (.CO(N1231), .S(N1230), .A(N426), .B(N472), .CI(N794));
ADDFXL inst_cellmath__63_0_I470 (.CO(N1233), .S(N1232), .A(N1215), .B(N748), .CI(N1226));
ADDFXL inst_cellmath__63_0_I471 (.CO(N1235), .S(N1234), .A(N1219), .B(N1217), .CI(N1228));
ADDFXL inst_cellmath__63_0_I472 (.CO(N1237), .S(N1236), .A(N1221), .B(N1230), .CI(N1232));
ADDFXL inst_cellmath__63_0_I473 (.CO(inst_cellmath__63_0_out1[9]), .S(inst_cellmath__63_0_out0[8]), .A(N1234), .B(N1223), .CI(N1236));
ADDHX1 inst_cellmath__63_0_I474 (.CO(N1241), .S(N1240), .A(N612), .B(N658));
ADDFX1 inst_cellmath__63_0_I475 (.CO(N1243), .S(N1242), .A(N704), .B(N750), .CI(N428));
ADDFX1 inst_cellmath__63_0_I476 (.CO(N1245), .S(N1244), .A(N474), .B(N520), .CI(N566));
ADDFX1 inst_cellmath__63_0_I477 (.CO(N1247), .S(N1246), .A(N796), .B(N842), .CI(N1227));
ADDFXL inst_cellmath__63_0_I478 (.CO(N1249), .S(N1248), .A(N1229), .B(N1240), .CI(N1231));
ADDFX1 inst_cellmath__63_0_I479 (.CO(N1251), .S(N1250), .A(N1244), .B(N1242), .CI(N1233));
ADDFXL inst_cellmath__63_0_I480 (.CO(N1253), .S(N1252), .A(N1235), .B(N1246), .CI(N1248));
ADDFXL inst_cellmath__63_0_I481 (.CO(inst_cellmath__63_0_out1[10]), .S(inst_cellmath__63_0_out0[9]), .A(N1250), .B(N1237), .CI(N1252));
ADDHX1 inst_cellmath__63_0_I482 (.CO(N1257), .S(N1256), .A(N660), .B(N430));
ADDFX1 inst_cellmath__63_0_I483 (.CO(N1259), .S(N1258), .A(N752), .B(N798), .CI(N476));
ADDFXL inst_cellmath__63_0_I484 (.CO(N1261), .S(N1260), .A(N522), .B(N568), .CI(N706));
ADDFX1 inst_cellmath__63_0_I485 (.CO(N1263), .S(N1262), .A(N890), .B(N614), .CI(N844));
ADDFX1 inst_cellmath__63_0_I486 (.CO(N1265), .S(N1264), .A(N1256), .B(N1241), .CI(N1243));
ADDFXL inst_cellmath__63_0_I487 (.CO(N1267), .S(N1266), .A(N1258), .B(N1245), .CI(N1260));
ADDFX1 inst_cellmath__63_0_I488 (.CO(N1269), .S(N1268), .A(N1262), .B(N1247), .CI(N1249));
ADDFXL inst_cellmath__63_0_I489 (.CO(N1271), .S(N1270), .A(N1251), .B(N1264), .CI(N1266));
ADDFXL inst_cellmath__63_0_I490 (.CO(inst_cellmath__63_0_out1[11]), .S(inst_cellmath__63_0_out0[10]), .A(N1253), .B(N1268), .CI(N1270));
ADDHX1 inst_cellmath__63_0_I491 (.CO(N1275), .S(N1274), .A(N708), .B(N478));
ADDFX1 inst_cellmath__63_0_I492 (.CO(N1277), .S(N1276), .A(N800), .B(N846), .CI(N524));
ADDFX1 inst_cellmath__63_0_I493 (.CO(N1279), .S(N1278), .A(N570), .B(N616), .CI(N754));
ADDFX1 inst_cellmath__63_0_I494 (.CO(N1281), .S(N1280), .A(N938), .B(N662), .CI(N892));
ADDFX1 inst_cellmath__63_0_I495 (.CO(N1283), .S(N1282), .A(N1257), .B(N432), .CI(N1274));
ADDFX1 inst_cellmath__63_0_I496 (.CO(N1285), .S(N1284), .A(N1261), .B(N1259), .CI(N1263));
ADDFX1 inst_cellmath__63_0_I497 (.CO(N1287), .S(N1286), .A(N1278), .B(N1276), .CI(N1280));
ADDFX1 inst_cellmath__63_0_I498 (.CO(N1289), .S(N1288), .A(N1282), .B(N1265), .CI(N1267));
ADDFX1 inst_cellmath__63_0_I499 (.CO(N1291), .S(N1290), .A(N1269), .B(N1284), .CI(N1286));
ADDFXL inst_cellmath__63_0_I500 (.CO(inst_cellmath__63_0_out1[12]), .S(inst_cellmath__63_0_out0[11]), .A(N1288), .B(N1271), .CI(N1290));
ADDHX1 inst_cellmath__63_0_I501 (.CO(N1295), .S(N1294), .A(N756), .B(N434));
ADDFX1 inst_cellmath__63_0_I502 (.CO(N1297), .S(N1296), .A(N848), .B(N894), .CI(N572));
ADDFX1 inst_cellmath__63_0_I503 (.CO(N1299), .S(N1298), .A(N618), .B(N664), .CI(N526));
ADDFX1 inst_cellmath__63_0_I504 (.CO(N1301), .S(N1300), .A(N802), .B(N710), .CI(N986));
ADDFX1 inst_cellmath__63_0_I505 (.CO(N1303), .S(N1302), .A(N940), .B(N480), .CI(N1275));
ADDFHX1 inst_cellmath__63_0_I506 (.CO(N1305), .S(N1304), .A(N1277), .B(N1294), .CI(N1279));
ADDFX1 inst_cellmath__63_0_I507 (.CO(N1307), .S(N1306), .A(N1296), .B(N1281), .CI(N1298));
ADDFX1 inst_cellmath__63_0_I508 (.CO(N1309), .S(N1308), .A(N1283), .B(N1300), .CI(N1302));
ADDFHX1 inst_cellmath__63_0_I509 (.CO(N1311), .S(N1310), .A(N1304), .B(N1285), .CI(N1287));
ADDFX1 inst_cellmath__63_0_I510 (.CO(N1313), .S(N1312), .A(N1289), .B(N1306), .CI(N1308));
ADDFXL inst_cellmath__63_0_I511 (.CO(inst_cellmath__63_0_out1[13]), .S(inst_cellmath__63_0_out0[12]), .A(N1310), .B(N1291), .CI(N1312));
ADDHX1 inst_cellmath__63_0_I512 (.CO(N1317), .S(N1316), .A(N804), .B(N482));
ADDFX1 inst_cellmath__63_0_I513 (.CO(N1319), .S(N1318), .A(N896), .B(N942), .CI(N620));
ADDFX1 inst_cellmath__63_0_I514 (.CO(N1321), .S(N1320), .A(N666), .B(N712), .CI(N574));
ADDFX1 inst_cellmath__63_0_I515 (.CO(N1323), .S(N1322), .A(N436), .B(N758), .CI(N850));
ADDFX1 inst_cellmath__63_0_I516 (.CO(N1325), .S(N1324), .A(N988), .B(N1034), .CI(N528));
ADDFXL inst_cellmath__63_0_I517 (.CO(N1327), .S(N1326), .A(N1316), .B(N1295), .CI(N1299));
ADDFX1 inst_cellmath__63_0_I518 (.CO(N1329), .S(N1328), .A(N1301), .B(N1297), .CI(N1318));
ADDFX1 inst_cellmath__63_0_I519 (.CO(N1331), .S(N1330), .A(N1322), .B(N1320), .CI(N1303));
ADDFXL inst_cellmath__63_0_I520 (.CO(N1333), .S(N1332), .A(N1305), .B(N1324), .CI(N1326));
ADDFX1 inst_cellmath__63_0_I521 (.CO(N1335), .S(N1334), .A(N1328), .B(N1307), .CI(N1309));
ADDFXL inst_cellmath__63_0_I522 (.CO(N1337), .S(N1336), .A(N1311), .B(N1330), .CI(N1332));
ADDFXL inst_cellmath__63_0_I523 (.CO(inst_cellmath__63_0_out1[14]), .S(inst_cellmath__63_0_out0[13]), .A(N1334), .B(N1313), .CI(N1336));
ADDHX1 inst_cellmath__63_0_I524 (.CO(N1341), .S(N1340), .A(N852), .B(N530));
ADDFX1 inst_cellmath__63_0_I525 (.CO(N1343), .S(N1342), .A(N438), .B(N990), .CI(N484));
ADDFX1 inst_cellmath__63_0_I526 (.CO(N1345), .S(N1344), .A(N760), .B(N944), .CI(N668));
ADDFX1 inst_cellmath__63_0_I527 (.CO(N1347), .S(N1346), .A(N806), .B(N714), .CI(N898));
ADDFX1 inst_cellmath__63_0_I528 (.CO(N1349), .S(N1348), .A(N1082), .B(N622), .CI(N1036));
ADDFX1 inst_cellmath__63_0_I529 (.CO(N1351), .S(N1350), .A(N1317), .B(N576), .CI(N1340));
ADDFX1 inst_cellmath__63_0_I530 (.CO(N1353), .S(N1352), .A(N1321), .B(N1319), .CI(N1323));
ADDFX1 inst_cellmath__63_0_I531 (.CO(N1355), .S(N1354), .A(N1342), .B(N1325), .CI(N1346));
ADDFX1 inst_cellmath__63_0_I532 (.CO(N1357), .S(N1356), .A(N1348), .B(N1344), .CI(N1327));
ADDFX1 inst_cellmath__63_0_I533 (.CO(N1359), .S(N1358), .A(N1329), .B(N1350), .CI(N1331));
ADDFX1 inst_cellmath__63_0_I534 (.CO(N1361), .S(N1360), .A(N1354), .B(N1352), .CI(N1333));
ADDFX1 inst_cellmath__63_0_I535 (.CO(N1363), .S(N1362), .A(N1335), .B(N1356), .CI(N1358));
ADDFX1 inst_cellmath__63_0_I536 (.CO(inst_cellmath__63_0_out1[15]), .S(inst_cellmath__63_0_out0[14]), .A(N1360), .B(N1337), .CI(N1362));
XNOR2X1 hap1_A_I716 (.Y(N1366), .A(N1130), .B(N992));
OR2XL hap1_A_I717 (.Y(N1367), .A(N1130), .B(N992));
ADDFX1 inst_cellmath__63_0_I538 (.CO(N1371), .S(N1370), .A(N486), .B(N900), .CI(N762));
ADDFXL inst_cellmath__63_0_I539 (.CO(N1373), .S(N1372), .A(N440), .B(N1038), .CI(N854));
ADDFX1 inst_cellmath__63_0_I540 (.CO(N1375), .S(N1374), .A(N532), .B(N808), .CI(N578));
ADDFXL inst_cellmath__63_0_I541 (.CO(N1377), .S(N1376), .A(N946), .B(N716), .CI(N670));
ADDFX1 inst_cellmath__63_0_I542 (.CO(N1379), .S(N1378), .A(N1084), .B(N624), .CI(N1341));
ADDFX1 inst_cellmath__63_0_I543 (.CO(N1381), .S(N1380), .A(N1343), .B(N1366), .CI(N1347));
ADDFX1 inst_cellmath__63_0_I544 (.CO(N1383), .S(N1382), .A(N1349), .B(N1345), .CI(N1372));
ADDFX1 inst_cellmath__63_0_I545 (.CO(N1385), .S(N1384), .A(N1374), .B(N1370), .CI(N1376));
ADDFX1 inst_cellmath__63_0_I546 (.CO(N1387), .S(N1386), .A(N1378), .B(N1351), .CI(N1353));
ADDFX1 inst_cellmath__63_0_I547 (.CO(N1389), .S(N1388), .A(N1380), .B(N1355), .CI(N1382));
ADDFX1 inst_cellmath__63_0_I548 (.CO(N1391), .S(N1390), .A(N1384), .B(N1357), .CI(N1359));
ADDFX1 inst_cellmath__63_0_I549 (.CO(N1393), .S(N1392), .A(N1361), .B(N1386), .CI(N1388));
ADDFX1 inst_cellmath__63_0_I550 (.CO(inst_cellmath__63_0_out1[16]), .S(inst_cellmath__63_0_out0[15]), .A(N1363), .B(N1390), .CI(N1392));
ADDFXL inst_cellmath__63_0_I551 (.CO(N1397), .S(N1396), .A(N1132), .B(N442), .CI(N856));
ADDFX1 inst_cellmath__63_0_I552 (.CO(N1399), .S(N1398), .A(N1040), .B(N948), .CI(N810));
ADDFXL inst_cellmath__63_0_I553 (.CO(N1401), .S(N1400), .A(N488), .B(N1086), .CI(N902));
ADDFXL inst_cellmath__63_0_I554 (.CO(N1403), .S(N1402), .A(N580), .B(N534), .CI(N626));
ADDFXL inst_cellmath__63_0_I555 (.CO(N1405), .S(N1404), .A(N994), .B(N764), .CI(N718));
ADDFXL inst_cellmath__63_0_I556 (.CO(N1407), .S(N1406), .A(N1367), .B(N672), .CI(N1373));
ADDFXL inst_cellmath__63_0_I557 (.CO(N1409), .S(N1408), .A(N1375), .B(N1371), .CI(N1377));
ADDFXL inst_cellmath__63_0_I558 (.CO(N1411), .S(N1410), .A(N1400), .B(N1396), .CI(N1402));
ADDFX1 inst_cellmath__63_0_I559 (.CO(N1413), .S(N1412), .A(N1404), .B(N1398), .CI(N1379));
ADDFXL inst_cellmath__63_0_I560 (.CO(N1415), .S(N1414), .A(N1406), .B(N1381), .CI(N1383));
ADDFXL inst_cellmath__63_0_I561 (.CO(N1417), .S(N1416), .A(N1408), .B(N1385), .CI(N1410));
ADDFXL inst_cellmath__63_0_I562 (.CO(N1419), .S(N1418), .A(N1387), .B(N1412), .CI(N1414));
ADDFX1 inst_cellmath__63_0_I563 (.CO(N1421), .S(N1420), .A(N1416), .B(N1389), .CI(N1391));
ADDFX1 inst_cellmath__63_0_I564 (.CO(inst_cellmath__63_0_out1[17]), .S(inst_cellmath__63_0_out0[16]), .A(N1393), .B(N1418), .CI(N1420));
ADDFXL inst_cellmath__63_0_I565 (.CO(N1425), .S(N1424), .A(N1134), .B(N444), .CI(N490));
ADDFXL inst_cellmath__63_0_I566 (.CO(N1427), .S(N1426), .A(N536), .B(N996), .CI(N950));
ADDFX1 inst_cellmath__63_0_I567 (.CO(N1429), .S(N1428), .A(N904), .B(N582), .CI(N812));
ADDFXL inst_cellmath__63_0_I568 (.CO(N1431), .S(N1430), .A(N858), .B(N1088), .CI(N766));
ADDFXL inst_cellmath__63_0_I569 (.CO(N1433), .S(N1432), .A(N1042), .B(N628), .CI(N674));
ADDFX1 inst_cellmath__63_0_I570 (.CO(N1435), .S(N1434), .A(N1397), .B(N720), .CI(N1399));
ADDFX1 inst_cellmath__63_0_I571 (.CO(N1437), .S(N1436), .A(N1401), .B(N1424), .CI(N1403));
ADDFXL inst_cellmath__63_0_I572 (.CO(N1439), .S(N1438), .A(N1426), .B(N1405), .CI(N1430));
ADDFX1 inst_cellmath__63_0_I573 (.CO(N1441), .S(N1440), .A(N1432), .B(N1428), .CI(N1407));
ADDFX1 inst_cellmath__63_0_I574 (.CO(N1443), .S(N1442), .A(N1434), .B(N1409), .CI(N1411));
ADDFXL inst_cellmath__63_0_I575 (.CO(N1445), .S(N1444), .A(N1413), .B(N1436), .CI(N1438));
ADDFXL inst_cellmath__63_0_I576 (.CO(N1447), .S(N1446), .A(N1415), .B(N1440), .CI(N1417));
ADDFXL inst_cellmath__63_0_I577 (.CO(N1449), .S(N1448), .A(N1444), .B(N1442), .CI(N1419));
ADDFXL inst_cellmath__63_0_I578 (.CO(inst_cellmath__63_0_out1[18]), .S(inst_cellmath__63_0_out0[17]), .A(N1421), .B(N1446), .CI(N1448));
INVXL fap1_A_I718 (.Y(N1803), .A(N1871));
ADDFX1 fap1_A_I719 (.CO(N1453), .S(N1452), .A(N1136), .B(N492), .CI(N1803));
ADDFXL inst_cellmath__63_0_I580 (.CO(N1457), .S(N1456), .A(N1044), .B(N538), .CI(N952));
ADDFXL inst_cellmath__63_0_I581 (.CO(N1459), .S(N1458), .A(N630), .B(N584), .CI(N906));
ADDFXL inst_cellmath__63_0_I582 (.CO(N1461), .S(N1460), .A(N860), .B(N998), .CI(N722));
ADDFX1 inst_cellmath__63_0_I583 (.CO(N1463), .S(N1462), .A(N1090), .B(N676), .CI(N814));
ADDFX1 inst_cellmath__63_0_I584 (.CO(N1465), .S(N1464), .A(N1425), .B(N768), .CI(N1427));
ADDFX1 inst_cellmath__63_0_I585 (.CO(N1467), .S(N1466), .A(N1431), .B(N1429), .CI(N1433));
ADDFXL inst_cellmath__63_0_I586 (.CO(N1469), .S(N1468), .A(N1456), .B(N1452), .CI(N1458));
ADDFX1 inst_cellmath__63_0_I587 (.CO(N1471), .S(N1470), .A(N1462), .B(N1460), .CI(N1435));
ADDFX1 inst_cellmath__63_0_I588 (.CO(N1473), .S(N1472), .A(N1464), .B(N1437), .CI(N1439));
ADDFX1 inst_cellmath__63_0_I589 (.CO(N1475), .S(N1474), .A(N1441), .B(N1466), .CI(N1468));
ADDFXL inst_cellmath__63_0_I590 (.CO(N1477), .S(N1476), .A(N1443), .B(N1470), .CI(N1445));
ADDFXL inst_cellmath__63_0_I591 (.CO(N1479), .S(N1478), .A(N1474), .B(N1472), .CI(N1447));
ADDFXL inst_cellmath__63_0_I592 (.CO(inst_cellmath__63_0_out1[19]), .S(inst_cellmath__63_0_out0[18]), .A(N1449), .B(N1476), .CI(N1478));
ADDFX1 inst_cellmath__63_0_I593 (.CO(N1483), .S(N1482), .A(N1871), .B(N1878), .CI(N540));
ADDFX1 inst_cellmath__63_0_I594 (.CO(N1485), .S(N1484), .A(N1092), .B(N586), .CI(N1138));
ADDFX1 inst_cellmath__63_0_I595 (.CO(N1487), .S(N1486), .A(N1000), .B(N632), .CI(N908));
ADDFX1 inst_cellmath__63_0_I596 (.CO(N1489), .S(N1488), .A(N954), .B(N678), .CI(N862));
ADDFX1 inst_cellmath__63_0_I597 (.CO(N1491), .S(N1490), .A(N1482), .B(N1046), .CI(N770));
ADDFXL inst_cellmath__63_0_I598 (.CO(N1493), .S(N1492), .A(N816), .B(N724), .CI(N1453));
ADDFXL inst_cellmath__63_0_I599 (.CO(N1495), .S(N1494), .A(N1459), .B(N1457), .CI(N1461));
ADDFX1 inst_cellmath__63_0_I600 (.CO(N1497), .S(N1496), .A(N1484), .B(N1463), .CI(N1486));
ADDFX1 inst_cellmath__63_0_I601 (.CO(N1499), .S(N1498), .A(N1488), .B(N1490), .CI(N1465));
ADDFXL inst_cellmath__63_0_I602 (.CO(N1501), .S(N1500), .A(N1467), .B(N1492), .CI(N1469));
ADDFXL inst_cellmath__63_0_I603 (.CO(N1503), .S(N1502), .A(N1471), .B(N1494), .CI(N1496));
ADDFXL inst_cellmath__63_0_I604 (.CO(N1505), .S(N1504), .A(N1473), .B(N1498), .CI(N1500));
ADDFXL inst_cellmath__63_0_I605 (.CO(N1507), .S(N1506), .A(N1502), .B(N1475), .CI(N1477));
ADDFXL inst_cellmath__63_0_I606 (.CO(inst_cellmath__63_0_out1[20]), .S(inst_cellmath__63_0_out0[19]), .A(N1479), .B(N1504), .CI(N1506));
ADDFXL inst_cellmath__63_0_I607 (.CO(N1511), .S(N1510), .A(N588), .B(N1885), .CI(N1140));
ADDFXL inst_cellmath__63_0_I608 (.CO(N1513), .S(N1512), .A(N1483), .B(N634), .CI(N680));
ADDFX1 inst_cellmath__63_0_I609 (.CO(N1515), .S(N1514), .A(N1048), .B(N726), .CI(N956));
ADDFX1 inst_cellmath__63_0_I610 (.CO(N1517), .S(N1516), .A(N772), .B(N1002), .CI(N910));
ADDFX1 inst_cellmath__63_0_I611 (.CO(N1519), .S(N1518), .A(N818), .B(N1094), .CI(N864));
ADDFXL inst_cellmath__63_0_I612 (.CO(N1521), .S(N1520), .A(N1510), .B(N1485), .CI(N1487));
ADDFX1 inst_cellmath__63_0_I613 (.CO(N1523), .S(N1522), .A(N1489), .B(N1491), .CI(N1512));
ADDFX1 inst_cellmath__63_0_I614 (.CO(N1525), .S(N1524), .A(N1514), .B(N1493), .CI(N1516));
ADDFXL inst_cellmath__63_0_I615 (.CO(N1527), .S(N1526), .A(N1495), .B(N1518), .CI(N1520));
ADDFX1 inst_cellmath__63_0_I616 (.CO(N1529), .S(N1528), .A(N1522), .B(N1497), .CI(N1499));
ADDFXL inst_cellmath__63_0_I617 (.CO(N1531), .S(N1530), .A(N1501), .B(N1524), .CI(N1526));
ADDFXL inst_cellmath__63_0_I618 (.CO(N1533), .S(N1532), .A(N1528), .B(N1503), .CI(N1505));
ADDFXL inst_cellmath__63_0_I619 (.CO(inst_cellmath__63_0_out1[21]), .S(inst_cellmath__63_0_out0[20]), .A(N1507), .B(N1530), .CI(N1532));
ADDFX1 inst_cellmath__63_0_I620 (.CO(N1537), .S(N1536), .A(N636), .B(N1892), .CI(N682));
ADDFX1 inst_cellmath__63_0_I621 (.CO(N1539), .S(N1538), .A(N728), .B(N1142), .CI(N1050));
ADDFX1 inst_cellmath__63_0_I622 (.CO(N1541), .S(N1540), .A(N1096), .B(N774), .CI(N1004));
ADDFX1 inst_cellmath__63_0_I623 (.CO(N1543), .S(N1542), .A(N958), .B(N820), .CI(N866));
ADDFX1 inst_cellmath__63_0_I624 (.CO(N1545), .S(N1544), .A(N1511), .B(N912), .CI(N1536));
ADDFX1 inst_cellmath__63_0_I625 (.CO(N1547), .S(N1546), .A(N1515), .B(N1513), .CI(N1517));
ADDFX1 inst_cellmath__63_0_I626 (.CO(N1549), .S(N1548), .A(N1538), .B(N1519), .CI(N1540));
ADDFXL inst_cellmath__63_0_I627 (.CO(N1551), .S(N1550), .A(N1521), .B(N1542), .CI(N1523));
ADDFX1 inst_cellmath__63_0_I628 (.CO(N1553), .S(N1552), .A(N1525), .B(N1544), .CI(N1546));
ADDFXL inst_cellmath__63_0_I629 (.CO(N1555), .S(N1554), .A(N1527), .B(N1548), .CI(N1550));
ADDFXL inst_cellmath__63_0_I630 (.CO(N1557), .S(N1556), .A(N1552), .B(N1529), .CI(N1531));
ADDFXL inst_cellmath__63_0_I631 (.CO(inst_cellmath__63_0_out1[22]), .S(inst_cellmath__63_0_out0[21]), .A(N1533), .B(N1554), .CI(N1556));
ADDFX1 inst_cellmath__63_0_I632 (.CO(N1561), .S(N1560), .A(N684), .B(N1899), .CI(N730));
ADDFX1 inst_cellmath__63_0_I633 (.CO(N1563), .S(N1562), .A(N776), .B(N1144), .CI(N1098));
ADDFX1 inst_cellmath__63_0_I634 (.CO(N1565), .S(N1564), .A(N868), .B(N822), .CI(N914));
ADDFX1 inst_cellmath__63_0_I635 (.CO(N1567), .S(N1566), .A(N1006), .B(N1052), .CI(N960));
ADDFX1 inst_cellmath__63_0_I636 (.CO(N1569), .S(N1568), .A(N1560), .B(N1537), .CI(N1539));
ADDFX1 inst_cellmath__63_0_I637 (.CO(N1571), .S(N1570), .A(N1543), .B(N1541), .CI(N1562));
ADDFX1 inst_cellmath__63_0_I638 (.CO(N1573), .S(N1572), .A(N1566), .B(N1564), .CI(N1545));
ADDFX1 inst_cellmath__63_0_I639 (.CO(N1575), .S(N1574), .A(N1568), .B(N1547), .CI(N1549));
ADDFX1 inst_cellmath__63_0_I640 (.CO(N1577), .S(N1576), .A(N1551), .B(N1570), .CI(N1572));
ADDFXL inst_cellmath__63_0_I641 (.CO(N1579), .S(N1578), .A(N1574), .B(N1553), .CI(N1555));
ADDFXL inst_cellmath__63_0_I642 (.CO(inst_cellmath__63_0_out1[23]), .S(inst_cellmath__63_0_out0[22]), .A(N1557), .B(N1576), .CI(N1578));
ADDFX1 inst_cellmath__63_0_I643 (.CO(N1583), .S(N1582), .A(N732), .B(N1906), .CI(N778));
ADDFX1 inst_cellmath__63_0_I644 (.CO(N1585), .S(N1584), .A(N824), .B(N1146), .CI(N870));
ADDFX1 inst_cellmath__63_0_I645 (.CO(N1587), .S(N1586), .A(N1100), .B(N916), .CI(N1054));
ADDFX1 inst_cellmath__63_0_I646 (.CO(N1589), .S(N1588), .A(N1008), .B(N962), .CI(N1561));
ADDFX1 inst_cellmath__63_0_I647 (.CO(N1591), .S(N1590), .A(N1563), .B(N1582), .CI(N1565));
ADDFX1 inst_cellmath__63_0_I648 (.CO(N1593), .S(N1592), .A(N1584), .B(N1567), .CI(N1586));
ADDFX1 inst_cellmath__63_0_I649 (.CO(N1595), .S(N1594), .A(N1569), .B(N1588), .CI(N1571));
ADDFX1 inst_cellmath__63_0_I650 (.CO(N1597), .S(N1596), .A(N1573), .B(N1590), .CI(N1592));
ADDFX1 inst_cellmath__63_0_I651 (.CO(N1599), .S(N1598), .A(N1594), .B(N1575), .CI(N1577));
ADDFX1 inst_cellmath__63_0_I652 (.CO(inst_cellmath__63_0_out1[24]), .S(inst_cellmath__63_0_out0[23]), .A(N1579), .B(N1596), .CI(N1598));
ADDFX1 inst_cellmath__63_0_I653 (.CO(N1603), .S(N1602), .A(N780), .B(N1913), .CI(N826));
ADDFX1 inst_cellmath__63_0_I654 (.CO(N1605), .S(N1604), .A(N872), .B(N1148), .CI(N918));
ADDFX1 inst_cellmath__63_0_I655 (.CO(N1607), .S(N1606), .A(N1102), .B(N964), .CI(N1010));
ADDFX1 inst_cellmath__63_0_I656 (.CO(N1609), .S(N1608), .A(N1583), .B(N1056), .CI(N1602));
ADDFX1 inst_cellmath__63_0_I657 (.CO(N1611), .S(N1610), .A(N1587), .B(N1585), .CI(N1589));
ADDFX1 inst_cellmath__63_0_I658 (.CO(N1613), .S(N1612), .A(N1606), .B(N1604), .CI(N1591));
ADDFX1 inst_cellmath__63_0_I659 (.CO(N1615), .S(N1614), .A(N1593), .B(N1608), .CI(N1610));
ADDFX1 inst_cellmath__63_0_I660 (.CO(N1617), .S(N1616), .A(N1612), .B(N1595), .CI(N1597));
ADDFX1 inst_cellmath__63_0_I661 (.CO(inst_cellmath__63_0_out1[25]), .S(inst_cellmath__63_0_out0[24]), .A(N1599), .B(N1614), .CI(N1616));
ADDFX1 inst_cellmath__63_0_I662 (.CO(N1621), .S(N1620), .A(N828), .B(N1920), .CI(N874));
ADDFX1 inst_cellmath__63_0_I663 (.CO(N1623), .S(N1622), .A(N920), .B(N1150), .CI(N966));
ADDFX1 inst_cellmath__63_0_I664 (.CO(N1625), .S(N1624), .A(N1058), .B(N1012), .CI(N1104));
ADDFX1 inst_cellmath__63_0_I665 (.CO(N1627), .S(N1626), .A(N1620), .B(N1603), .CI(N1605));
ADDFX1 inst_cellmath__63_0_I666 (.CO(N1629), .S(N1628), .A(N1622), .B(N1607), .CI(N1609));
ADDFX1 inst_cellmath__63_0_I667 (.CO(N1631), .S(N1630), .A(N1611), .B(N1624), .CI(N1626));
ADDFX1 inst_cellmath__63_0_I668 (.CO(N1633), .S(N1632), .A(N1628), .B(N1613), .CI(N1615));
ADDFX1 inst_cellmath__63_0_I669 (.CO(inst_cellmath__63_0_out1[26]), .S(inst_cellmath__63_0_out0[25]), .A(N1617), .B(N1630), .CI(N1632));
ADDFX1 inst_cellmath__63_0_I670 (.CO(N1637), .S(N1636), .A(N876), .B(N1921), .CI(N922));
ADDFX1 inst_cellmath__63_0_I671 (.CO(N1639), .S(N1638), .A(N968), .B(N1152), .CI(N1014));
ADDFX1 inst_cellmath__63_0_I672 (.CO(N1641), .S(N1640), .A(N1106), .B(N1060), .CI(N1621));
ADDFX1 inst_cellmath__63_0_I673 (.CO(N1643), .S(N1642), .A(N1623), .B(N1636), .CI(N1625));
ADDFX1 inst_cellmath__63_0_I674 (.CO(N1645), .S(N1644), .A(N1640), .B(N1638), .CI(N1627));
ADDFX1 inst_cellmath__63_0_I675 (.CO(N1647), .S(N1646), .A(N1629), .B(N1642), .CI(N1644));
ADDFX1 inst_cellmath__63_0_I676 (.CO(inst_cellmath__63_0_out1[27]), .S(inst_cellmath__63_0_out0[26]), .A(N1633), .B(N1631), .CI(N1646));
ADDFX1 inst_cellmath__63_0_I677 (.CO(N1651), .S(N1650), .A(N924), .B(N1922), .CI(N970));
ADDFX1 inst_cellmath__63_0_I678 (.CO(N1653), .S(N1652), .A(N1016), .B(N1154), .CI(N1062));
ADDFX1 inst_cellmath__63_0_I679 (.CO(N1655), .S(N1654), .A(N1637), .B(N1108), .CI(N1650));
ADDFX1 inst_cellmath__63_0_I680 (.CO(N1657), .S(N1656), .A(N1641), .B(N1639), .CI(N1652));
ADDFX1 inst_cellmath__63_0_I681 (.CO(N1659), .S(N1658), .A(N1654), .B(N1643), .CI(N1645));
ADDFX1 inst_cellmath__63_0_I682 (.CO(inst_cellmath__63_0_out1[28]), .S(inst_cellmath__63_0_out0[27]), .A(N1647), .B(N1656), .CI(N1658));
ADDFX1 inst_cellmath__63_0_I683 (.CO(N1663), .S(N1662), .A(N972), .B(N1929), .CI(N1018));
ADDFX1 inst_cellmath__63_0_I684 (.CO(N1665), .S(N1664), .A(N1064), .B(N1156), .CI(N1110));
ADDFX1 inst_cellmath__63_0_I685 (.CO(N1667), .S(N1666), .A(N1662), .B(N1651), .CI(N1653));
ADDFX1 inst_cellmath__63_0_I686 (.CO(N1669), .S(N1668), .A(N1655), .B(N1664), .CI(N1666));
ADDFX1 inst_cellmath__63_0_I687 (.CO(inst_cellmath__63_0_out0[29]), .S(inst_cellmath__63_0_out0[28]), .A(N1659), .B(N1657), .CI(N1668));
ADDFX1 inst_cellmath__63_0_I688 (.CO(N1673), .S(N1672), .A(N1020), .B(N1930), .CI(N1158));
ADDFX1 inst_cellmath__63_0_I689 (.CO(N1675), .S(N1674), .A(N1112), .B(N1066), .CI(N1663));
ADDFX1 inst_cellmath__63_0_I690 (.CO(N1677), .S(N1676), .A(N1665), .B(N1672), .CI(N1674));
ADDFX1 inst_cellmath__63_0_I691 (.CO(inst_cellmath__63_0_out0[30]), .S(inst_cellmath__63_0_out1[29]), .A(N1676), .B(N1667), .CI(N1669));
ADDFX1 inst_cellmath__63_0_I692 (.CO(N1681), .S(N1680), .A(N1068), .B(N1931), .CI(N1160));
ADDFX1 inst_cellmath__63_0_I693 (.CO(N1683), .S(N1682), .A(N1673), .B(N1114), .CI(N1680));
ADDFX1 inst_cellmath__63_0_I694 (.CO(inst_cellmath__63_0_out0[31]), .S(inst_cellmath__63_0_out1[30]), .A(N1682), .B(N1675), .CI(N1677));
ADDFX1 inst_cellmath__63_0_I695 (.CO(N1687), .S(N1686), .A(N1116), .B(N1938), .CI(N1162));
ADDFX1 inst_cellmath__63_0_I696 (.CO(inst_cellmath__63_0_out0[32]), .S(inst_cellmath__63_0_out1[31]), .A(N1686), .B(N1681), .CI(N1683));
ADDFX1 inst_cellmath__63_0_I697 (.CO(inst_cellmath__63_0_out0[33]), .S(inst_cellmath__63_0_out1[32]), .A(N1164), .B(N1939), .CI(N1687));
assign inst_cellmath__63_0_out0[0] = 1'B0;
assign inst_cellmath__63_0_out0[34] = 1'B0;
assign inst_cellmath__63_0_out0[35] = 1'B0;
assign inst_cellmath__63_0_out0[36] = 1'B0;
assign inst_cellmath__63_0_out0[37] = 1'B0;
assign inst_cellmath__63_0_out0[38] = 1'B0;
assign inst_cellmath__63_0_out0[39] = 1'B0;
assign inst_cellmath__63_0_out1[34] = 1'B1;
assign inst_cellmath__63_0_out1[35] = 1'B1;
assign inst_cellmath__63_0_out1[36] = 1'B1;
assign inst_cellmath__63_0_out1[37] = 1'B1;
assign inst_cellmath__63_0_out1[38] = 1'B1;
assign inst_cellmath__63_0_out1[39] = 1'B1;
endmodule

module cynw_cm_float_rcp_inst_cellmath__64_0_bdw1471647203_bdw (
	inst_cellmath__64_0_out0,
	inst_cellmath__64_0_in0,
	inst_cellmath__64_0_in1,
	inst_cellmath__64_0_in2,
	inst_cellmath__64_0_in3,
	inst_cellmath__64_0_in4
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__64_0_out0;
input [52:28] inst_cellmath__64_0_in0;
input [39:0] inst_cellmath__64_0_in1,
	inst_cellmath__64_0_in2,
	inst_cellmath__64_0_in3,
	inst_cellmath__64_0_in4;
wire N1509,N1510,N1511,N1512,N1513,N1514,N1515 
	,N1516,N1517,N1518,N1519,N1520,N1521,N1522,N1523 
	,N1524,N1525,N1526,N1527,N1528,N1529,N1530,N1531 
	,N1532,N1533,N1534,N1535,N1536,N1537,N1538,N1539 
	,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547 
	,N1548,N1549,N1550,N1551,N1552,N1553,N1554,N1555 
	,N1556,N1557,N1558,N1559,N1560,N1561,N1562,N1563 
	,N1564,N1565,N1566,N1567,N1568,N1569,N1570,N1571 
	,N1572,N1573,N1574,N1577,N1578,N1579,N1580,N1581 
	,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589 
	,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597 
	,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605 
	,N1606,N1607,N1608,N1609,N1610,N1611,N1612,N1613 
	,N1614,N1615,N1616,N1617,N1618,N1619,N1620,N1621 
	,N1622,N1623,N1624,N1625,N1626,N1627,N1628,N1629 
	,N1630,N1631,N1632,N1633,N1634,N1635,N1636,N1637 
	,N1638,N1639,N1640,N1641,N1642,N1643,N1644,N1645 
	,N1646,N1647,N1648,N1649,N1650,N1651,N1652,N1653 
	,N1654,N1655,N1656,N1657,N1658,N1659,N1660,N1661 
	,N1662,N1663,N1664,N1665,N1666,N1667,N1668,N1669 
	,N1670,N1671,N1672,N1673,N1674,N1675,N1676,N1677 
	,N1678,N1679,N1680,N1681,N1682,N1683,N1684,N1685 
	,N1686,N1687,N1688,N1689,N1690,N1691,N1692,N1693 
	,N1694,N1695,N1696,N1697,N1698,N1699,N1700,N1701 
	,N1702,N1703,N1704,N1705,N1706,N1707,N1708,N1709 
	,N1710,N1711,N1712,N1713,N1714,N1715,N1716,N1717 
	,N1718,N1719,N1720,N1721,N1722,N1723,N1724,N1725 
	,N1726,N1727,N1728,N1729,N1730,N1731,N1732,N1733 
	,N1734,N1735,N1736,N1737,N1738,N1739,N1740,N1741 
	,N1742,N1743,N1744,N1745,N1746,N1747,N1748,N1749 
	,N1750,N1751,N1752,N1753,N1754,N1755,N1756,N1757 
	,N1759,N1760,N1761,N1762,N1763,N1764,N1765,N1767 
	,N1768,N1769,N1770,N1771,N1772,N1773,N1774,N1775 
	,N1776,N1777,N1778,N1779,N1780,N1781,N1782,N1783 
	,N1784,N1785,N1786,N1787,N1788,N1789,N1790,N1791 
	,N1792,N1793,N1794,N1795,N1796,N1799,N1807,N1815 
	,N1827,N1839,N1855,N1871,N1891,N1911,N1935,N1959 
	,N1987,N2015,N2047,N2079,N2102,N2105,N2108,N2111 
	,N2114,N2117,N2120,N2123,N2126,N2129,N2132,N2135 
	,N2138,N2141,N2144,N2161,N2163,N2164,N2165,N2166 
	,N2167,N2168,N2169,N2170,N2171,N2172,N2173,N2174 
	,N2175,N2176,N2177,N2178,N2179,N2180,N2181,N2182 
	,N2183,N2184,N2185,N2186,N2187,N2188,N2189,N2190 
	,N2191,N2192,N2193,N2194,N2195,N2196,N2197,N2198 
	,N2199,N2200,N2201,N2202,N2203,N2204,N2205,N2206 
	,N2207,N2208,N2209,N2210,N2215,N2219,N2223,N2231 
	,N2235,N2236,N2239,N2240,N2247,N2248,N2251,N2252 
	,N2255,N2256,N2263,N2264,N2267,N2268,N2271,N2272 
	,N2279,N2280,N2283,N2284,N2319,N2321,N2322,N2323 
	,N2324,N2325,N2326,N2327,N2328,N2329,N2330,N2331 
	,N2332,N2337,N2339,N2341,N2342,N2343,N2344,N2345 
	,N2346,N2347,N2348,N2357,N2359,N2361,N2363,N2432 
	,N2435,N2438,N2441,N2444,N2447,N2450,N2453,N2456 
	,N2459,N2462,N2471,N2474,N2483,N2486,N2495,N2498 
	,N2515,N2516,N2518,N2519,N2521,N2522,N2524,N2525 
	,N2527,N2528,N2530,N2531,N2533,N2534,N2536,N2537 
	,N2539,N2540,N2542,N2543,N2545,N2546,N2548,N2549 
	,N2551,N2552,N2554,N2555,N2557,N2558,N2560,N2561 
	,N2606,N2678,N2680,N2689,N2691,N2707,N2709,N2718 
	,N2720,N2736,N2738,N2747,N2749,N2765,N2767,N2776 
	,N2778,N2875,N2876,N2882,N2883,N2893,N2894,N2908 
	,N2909,N2927,N2928,N2950,N2951,N2977,N2978,N3020 
	,N3028,N3036,N3044,N3050,N3053,N3054,N3057,N3060 
	,N3063,N3066,N3069,N3072,N3073,N3074,N3075,N3076 
	,N3077,N3078,N3079,N3093,N3099,N3105,N3111,N3114 
	,N3121,N3128,N3135;
ADDHX1 inst_cellmath__64_0_I412 (.CO(N1510), .S(N1509), .A(inst_cellmath__64_0_in1[0]), .B(inst_cellmath__64_0_in4[0]));
ADDHX1 inst_cellmath__64_0_I413 (.CO(N1512), .S(N1511), .A(inst_cellmath__64_0_in4[1]), .B(inst_cellmath__64_0_in3[1]));
ADDFX1 inst_cellmath__64_0_I414 (.CO(N1514), .S(N1513), .A(N1511), .B(N1510), .CI(inst_cellmath__64_0_in2[1]));
ADDFX1 inst_cellmath__64_0_I415 (.CO(N1516), .S(N1515), .A(inst_cellmath__64_0_in3[2]), .B(inst_cellmath__64_0_in4[2]), .CI(N1512));
ADDFX1 inst_cellmath__64_0_I416 (.CO(N1518), .S(N1517), .A(inst_cellmath__64_0_in2[2]), .B(N1515), .CI(N1514));
ADDFX1 inst_cellmath__64_0_I417 (.CO(N1520), .S(N1519), .A(inst_cellmath__64_0_in3[3]), .B(inst_cellmath__64_0_in4[3]), .CI(N1516));
ADDFX1 inst_cellmath__64_0_I418 (.CO(N1522), .S(N1521), .A(inst_cellmath__64_0_in2[3]), .B(N1519), .CI(N1518));
ADDFX1 inst_cellmath__64_0_I419 (.CO(N1524), .S(N1523), .A(N1520), .B(inst_cellmath__64_0_in3[4]), .CI(inst_cellmath__64_0_in2[4]));
ADDFX1 inst_cellmath__64_0_I420 (.CO(N1526), .S(N1525), .A(inst_cellmath__64_0_in4[4]), .B(N1522), .CI(N1523));
ADDFX1 inst_cellmath__64_0_I421 (.CO(N1528), .S(N1527), .A(inst_cellmath__64_0_in3[5]), .B(N1524), .CI(inst_cellmath__64_0_in4[5]));
ADDFX1 inst_cellmath__64_0_I422 (.CO(N1530), .S(N1529), .A(N1526), .B(inst_cellmath__64_0_in2[5]), .CI(inst_cellmath__64_0_in1[5]));
ADDFX1 inst_cellmath__64_0_I423 (.CO(N1532), .S(N1531), .A(inst_cellmath__64_0_in2[6]), .B(inst_cellmath__64_0_in4[6]), .CI(N1528));
ADDFX1 inst_cellmath__64_0_I424 (.CO(N1534), .S(N1533), .A(inst_cellmath__64_0_in1[6]), .B(inst_cellmath__64_0_in3[6]), .CI(N1530));
ADDFX1 inst_cellmath__64_0_I425 (.CO(N1536), .S(N1535), .A(inst_cellmath__64_0_in2[7]), .B(inst_cellmath__64_0_in4[7]), .CI(N1532));
ADDFX1 inst_cellmath__64_0_I426 (.CO(N1538), .S(N1537), .A(inst_cellmath__64_0_in3[7]), .B(inst_cellmath__64_0_in1[7]), .CI(N1534));
ADDFX1 inst_cellmath__64_0_I427 (.CO(N1540), .S(N1539), .A(inst_cellmath__64_0_in4[8]), .B(inst_cellmath__64_0_in2[8]), .CI(N1536));
ADDFX1 inst_cellmath__64_0_I428 (.CO(N1542), .S(N1541), .A(inst_cellmath__64_0_in3[8]), .B(inst_cellmath__64_0_in1[8]), .CI(N1538));
ADDFX1 inst_cellmath__64_0_I429 (.CO(N1544), .S(N1543), .A(inst_cellmath__64_0_in4[9]), .B(inst_cellmath__64_0_in2[9]), .CI(inst_cellmath__64_0_in1[9]));
ADDFX1 inst_cellmath__64_0_I430 (.CO(N1546), .S(N1545), .A(inst_cellmath__64_0_in3[9]), .B(N1540), .CI(N1543));
ADDFX1 inst_cellmath__64_0_I431 (.CO(N1548), .S(N1547), .A(inst_cellmath__64_0_in1[10]), .B(inst_cellmath__64_0_in2[10]), .CI(inst_cellmath__64_0_in4[10]));
ADDFX1 inst_cellmath__64_0_I432 (.CO(N1550), .S(N1549), .A(N1547), .B(N1544), .CI(inst_cellmath__64_0_in3[10]));
ADDFX1 inst_cellmath__64_0_I433 (.CO(N1552), .S(N1551), .A(inst_cellmath__64_0_in1[11]), .B(inst_cellmath__64_0_in2[11]), .CI(N1548));
ADDFHXL inst_cellmath__64_0_I434 (.CO(N1554), .S(N1553), .A(inst_cellmath__64_0_in3[11]), .B(inst_cellmath__64_0_in4[11]), .CI(N1551));
ADDFX1 inst_cellmath__64_0_I435 (.CO(N1556), .S(N1555), .A(inst_cellmath__64_0_in1[12]), .B(inst_cellmath__64_0_in2[12]), .CI(inst_cellmath__64_0_in4[12]));
ADDFX1 inst_cellmath__64_0_I436 (.CO(N1558), .S(N1557), .A(inst_cellmath__64_0_in3[12]), .B(N1552), .CI(N1555));
ADDFX1 inst_cellmath__64_0_I437 (.CO(N1560), .S(N1559), .A(inst_cellmath__64_0_in1[13]), .B(inst_cellmath__64_0_in2[13]), .CI(inst_cellmath__64_0_in4[13]));
ADDFX1 inst_cellmath__64_0_I438 (.CO(N1562), .S(N1561), .A(inst_cellmath__64_0_in3[13]), .B(N1556), .CI(N1559));
ADDFX1 inst_cellmath__64_0_I439 (.CO(N1564), .S(N1563), .A(inst_cellmath__64_0_in1[14]), .B(inst_cellmath__64_0_in2[14]), .CI(inst_cellmath__64_0_in4[14]));
ADDFX1 inst_cellmath__64_0_I440 (.CO(N1566), .S(N1565), .A(inst_cellmath__64_0_in3[14]), .B(N1560), .CI(N1563));
ADDHX1 inst_cellmath__64_0_I441 (.CO(N1568), .S(N1567), .A(inst_cellmath__64_0_in0[28]), .B(inst_cellmath__64_0_in2[15]));
ADDFX1 inst_cellmath__64_0_I442 (.CO(N1570), .S(N1569), .A(inst_cellmath__64_0_in1[15]), .B(N1567), .CI(inst_cellmath__64_0_in4[15]));
ADDFX1 inst_cellmath__64_0_I443 (.CO(N1572), .S(N1571), .A(inst_cellmath__64_0_in3[15]), .B(N1564), .CI(N1569));
INVXL fap1_A_I1339 (.Y(N2606), .A(inst_cellmath__64_0_in0[29]));
ADDFX1 fap1_A_I1340 (.CO(N1574), .S(N1573), .A(inst_cellmath__64_0_in2[16]), .B(N1568), .CI(N2606));
ADDFXL inst_cellmath__64_0_I445 (.CO(N1578), .S(N1577), .A(N1573), .B(inst_cellmath__64_0_in1[16]), .CI(inst_cellmath__64_0_in4[16]));
ADDFX1 inst_cellmath__64_0_I446 (.CO(N1580), .S(N1579), .A(inst_cellmath__64_0_in3[16]), .B(N1570), .CI(N1577));
ADDHX1 inst_cellmath__64_0_I447 (.CO(N1582), .S(N1581), .A(inst_cellmath__64_0_in0[29]), .B(inst_cellmath__64_0_in0[30]));
ADDFX1 inst_cellmath__64_0_I448 (.CO(N1584), .S(N1583), .A(inst_cellmath__64_0_in2[17]), .B(N1581), .CI(inst_cellmath__64_0_in1[17]));
ADDFXL inst_cellmath__64_0_I449 (.CO(N1586), .S(N1585), .A(inst_cellmath__64_0_in4[17]), .B(N1574), .CI(inst_cellmath__64_0_in3[17]));
ADDFX1 inst_cellmath__64_0_I450 (.CO(N1588), .S(N1587), .A(N1578), .B(N1583), .CI(N1585));
ADDHX1 inst_cellmath__64_0_I451 (.CO(N1590), .S(N1589), .A(inst_cellmath__64_0_in0[31]), .B(N1582));
ADDFX1 inst_cellmath__64_0_I452 (.CO(N1592), .S(N1591), .A(inst_cellmath__64_0_in2[18]), .B(N1589), .CI(inst_cellmath__64_0_in1[18]));
ADDFX1 inst_cellmath__64_0_I453 (.CO(N1594), .S(N1593), .A(N1584), .B(inst_cellmath__64_0_in4[18]), .CI(inst_cellmath__64_0_in3[18]));
ADDFX1 inst_cellmath__64_0_I454 (.CO(N1596), .S(N1595), .A(N1586), .B(N1591), .CI(N1593));
ADDHX1 inst_cellmath__64_0_I455 (.CO(N1598), .S(N1597), .A(inst_cellmath__64_0_in0[32]), .B(N1590));
ADDFX1 inst_cellmath__64_0_I456 (.CO(N1600), .S(N1599), .A(inst_cellmath__64_0_in2[19]), .B(N1597), .CI(inst_cellmath__64_0_in1[19]));
ADDFX1 inst_cellmath__64_0_I457 (.CO(N1602), .S(N1601), .A(N1592), .B(inst_cellmath__64_0_in4[19]), .CI(inst_cellmath__64_0_in3[19]));
ADDFXL inst_cellmath__64_0_I458 (.CO(N1604), .S(N1603), .A(N1594), .B(N1599), .CI(N1601));
ADDHX1 inst_cellmath__64_0_I459 (.CO(N1606), .S(N1605), .A(inst_cellmath__64_0_in0[33]), .B(N1598));
ADDFX1 inst_cellmath__64_0_I460 (.CO(N1608), .S(N1607), .A(inst_cellmath__64_0_in2[20]), .B(N1605), .CI(inst_cellmath__64_0_in1[20]));
ADDFX1 inst_cellmath__64_0_I461 (.CO(N1610), .S(N1609), .A(N1600), .B(inst_cellmath__64_0_in4[20]), .CI(inst_cellmath__64_0_in3[20]));
ADDFX1 inst_cellmath__64_0_I462 (.CO(N1612), .S(N1611), .A(N1602), .B(N1607), .CI(N1609));
ADDHX1 inst_cellmath__64_0_I463 (.CO(N1614), .S(N1613), .A(inst_cellmath__64_0_in0[34]), .B(N1606));
ADDFX1 inst_cellmath__64_0_I464 (.CO(N1616), .S(N1615), .A(inst_cellmath__64_0_in2[21]), .B(N1613), .CI(inst_cellmath__64_0_in1[21]));
ADDFX1 inst_cellmath__64_0_I465 (.CO(N1618), .S(N1617), .A(inst_cellmath__64_0_in3[21]), .B(inst_cellmath__64_0_in4[21]), .CI(N1608));
ADDFX1 inst_cellmath__64_0_I466 (.CO(N1620), .S(N1619), .A(N1610), .B(N1615), .CI(N1617));
ADDHX1 inst_cellmath__64_0_I467 (.CO(N1622), .S(N1621), .A(inst_cellmath__64_0_in0[35]), .B(N1614));
ADDFX1 inst_cellmath__64_0_I468 (.CO(N1624), .S(N1623), .A(inst_cellmath__64_0_in2[22]), .B(N1621), .CI(inst_cellmath__64_0_in4[22]));
ADDFX1 inst_cellmath__64_0_I469 (.CO(N1626), .S(N1625), .A(inst_cellmath__64_0_in1[22]), .B(inst_cellmath__64_0_in3[22]), .CI(N1623));
ADDFX1 inst_cellmath__64_0_I470 (.CO(N1628), .S(N1627), .A(N1618), .B(N1616), .CI(N1625));
ADDHX1 inst_cellmath__64_0_I471 (.CO(N1630), .S(N1629), .A(inst_cellmath__64_0_in0[36]), .B(N1622));
ADDFX1 inst_cellmath__64_0_I472 (.CO(N1632), .S(N1631), .A(inst_cellmath__64_0_in4[23]), .B(N1629), .CI(inst_cellmath__64_0_in3[23]));
ADDFX1 inst_cellmath__64_0_I473 (.CO(N1634), .S(N1633), .A(inst_cellmath__64_0_in1[23]), .B(inst_cellmath__64_0_in2[23]), .CI(N1631));
ADDFX1 inst_cellmath__64_0_I474 (.CO(N1636), .S(N1635), .A(N1633), .B(N1624), .CI(N1626));
ADDHX1 inst_cellmath__64_0_I475 (.CO(N1638), .S(N1637), .A(inst_cellmath__64_0_in0[37]), .B(N1630));
ADDFX1 inst_cellmath__64_0_I476 (.CO(N1640), .S(N1639), .A(inst_cellmath__64_0_in4[24]), .B(N1637), .CI(inst_cellmath__64_0_in3[24]));
ADDFX1 inst_cellmath__64_0_I477 (.CO(N1642), .S(N1641), .A(inst_cellmath__64_0_in2[24]), .B(N1639), .CI(inst_cellmath__64_0_in1[24]));
ADDFX1 inst_cellmath__64_0_I478 (.CO(N1644), .S(N1643), .A(N1641), .B(N1632), .CI(N1634));
ADDHX1 inst_cellmath__64_0_I479 (.CO(N1646), .S(N1645), .A(inst_cellmath__64_0_in4[25]), .B(inst_cellmath__64_0_in3[25]));
ADDFX1 inst_cellmath__64_0_I480 (.CO(N1648), .S(N1647), .A(inst_cellmath__64_0_in0[38]), .B(N1645), .CI(N1638));
ADDFX1 inst_cellmath__64_0_I481 (.CO(N1650), .S(N1649), .A(N1640), .B(N1647), .CI(inst_cellmath__64_0_in2[25]));
ADDFX1 inst_cellmath__64_0_I482 (.CO(N1652), .S(N1651), .A(N1649), .B(inst_cellmath__64_0_in1[25]), .CI(N1642));
ADDHX1 inst_cellmath__64_0_I483 (.CO(N1654), .S(N1653), .A(inst_cellmath__64_0_in4[26]), .B(inst_cellmath__64_0_in3[26]));
ADDFX1 inst_cellmath__64_0_I484 (.CO(N1656), .S(N1655), .A(N1653), .B(N1646), .CI(inst_cellmath__64_0_in0[39]));
ADDFX1 inst_cellmath__64_0_I485 (.CO(N1658), .S(N1657), .A(N1648), .B(N1655), .CI(inst_cellmath__64_0_in2[26]));
ADDFX1 inst_cellmath__64_0_I486 (.CO(N1660), .S(N1659), .A(N1650), .B(inst_cellmath__64_0_in1[26]), .CI(N1657));
ADDHX1 inst_cellmath__64_0_I487 (.CO(N1662), .S(N1661), .A(inst_cellmath__64_0_in4[27]), .B(inst_cellmath__64_0_in3[27]));
ADDFX1 inst_cellmath__64_0_I488 (.CO(N1664), .S(N1663), .A(N1661), .B(N1654), .CI(inst_cellmath__64_0_in0[40]));
ADDFX1 inst_cellmath__64_0_I489 (.CO(N1666), .S(N1665), .A(N1663), .B(N1656), .CI(inst_cellmath__64_0_in1[27]));
ADDFX1 inst_cellmath__64_0_I490 (.CO(N1668), .S(N1667), .A(N1658), .B(inst_cellmath__64_0_in2[27]), .CI(N1665));
ADDHX1 inst_cellmath__64_0_I491 (.CO(N1670), .S(N1669), .A(inst_cellmath__64_0_in4[28]), .B(inst_cellmath__64_0_in3[28]));
ADDFX1 inst_cellmath__64_0_I492 (.CO(N1672), .S(N1671), .A(N1669), .B(N1662), .CI(inst_cellmath__64_0_in0[41]));
ADDFX1 inst_cellmath__64_0_I493 (.CO(N1674), .S(N1673), .A(N1671), .B(N1664), .CI(inst_cellmath__64_0_in2[28]));
ADDFX1 inst_cellmath__64_0_I494 (.CO(N1676), .S(N1675), .A(N1673), .B(inst_cellmath__64_0_in1[28]), .CI(N1666));
ADDHX1 inst_cellmath__64_0_I495 (.CO(N1678), .S(N1677), .A(inst_cellmath__64_0_in4[29]), .B(inst_cellmath__64_0_in3[29]));
ADDFX1 inst_cellmath__64_0_I496 (.CO(N1680), .S(N1679), .A(N1677), .B(N1670), .CI(inst_cellmath__64_0_in0[42]));
ADDFX1 inst_cellmath__64_0_I497 (.CO(N1682), .S(N1681), .A(N1679), .B(N1672), .CI(inst_cellmath__64_0_in2[29]));
ADDFX1 inst_cellmath__64_0_I498 (.CO(N1684), .S(N1683), .A(N1681), .B(inst_cellmath__64_0_in1[29]), .CI(N1674));
ADDHX1 inst_cellmath__64_0_I499 (.CO(N1686), .S(N1685), .A(inst_cellmath__64_0_in4[30]), .B(inst_cellmath__64_0_in3[30]));
ADDFX1 inst_cellmath__64_0_I500 (.CO(N1688), .S(N1687), .A(N1685), .B(N1678), .CI(inst_cellmath__64_0_in0[43]));
ADDFX1 inst_cellmath__64_0_I501 (.CO(N1690), .S(N1689), .A(N1687), .B(N1680), .CI(inst_cellmath__64_0_in2[30]));
ADDFX1 inst_cellmath__64_0_I502 (.CO(N1692), .S(N1691), .A(N1689), .B(inst_cellmath__64_0_in1[30]), .CI(N1682));
ADDHX1 inst_cellmath__64_0_I503 (.CO(N1694), .S(N1693), .A(inst_cellmath__64_0_in4[31]), .B(inst_cellmath__64_0_in3[31]));
ADDFX1 inst_cellmath__64_0_I504 (.CO(N1696), .S(N1695), .A(N1693), .B(N1686), .CI(inst_cellmath__64_0_in0[44]));
ADDFX1 inst_cellmath__64_0_I505 (.CO(N1698), .S(N1697), .A(N1695), .B(N1688), .CI(inst_cellmath__64_0_in2[31]));
ADDFX1 inst_cellmath__64_0_I506 (.CO(N1700), .S(N1699), .A(N1697), .B(inst_cellmath__64_0_in1[31]), .CI(N1690));
ADDHX1 inst_cellmath__64_0_I507 (.CO(N1702), .S(N1701), .A(inst_cellmath__64_0_in4[32]), .B(inst_cellmath__64_0_in3[32]));
ADDFX1 inst_cellmath__64_0_I508 (.CO(N1704), .S(N1703), .A(N1701), .B(N1694), .CI(inst_cellmath__64_0_in0[45]));
ADDFX1 inst_cellmath__64_0_I509 (.CO(N1706), .S(N1705), .A(N1703), .B(N1696), .CI(inst_cellmath__64_0_in2[32]));
ADDFX1 inst_cellmath__64_0_I510 (.CO(N1708), .S(N1707), .A(inst_cellmath__64_0_in1[32]), .B(N1705), .CI(N1698));
ADDHX1 inst_cellmath__64_0_I511 (.CO(N1710), .S(N1709), .A(inst_cellmath__64_0_in4[33]), .B(inst_cellmath__64_0_in3[33]));
ADDFX1 inst_cellmath__64_0_I512 (.CO(N1712), .S(N1711), .A(N1709), .B(N1702), .CI(inst_cellmath__64_0_in2[33]));
ADDFX1 inst_cellmath__64_0_I513 (.CO(N1714), .S(N1713), .A(inst_cellmath__64_0_in0[46]), .B(N1711), .CI(N1704));
ADDFX1 inst_cellmath__64_0_I514 (.CO(N1716), .S(N1715), .A(N1713), .B(inst_cellmath__64_0_in1[33]), .CI(N1706));
ADDHX1 inst_cellmath__64_0_I515 (.CO(N1718), .S(N1717), .A(inst_cellmath__64_0_in2[34]), .B(inst_cellmath__64_0_in1[34]));
ADDFX1 inst_cellmath__64_0_I516 (.CO(N1720), .S(N1719), .A(inst_cellmath__64_0_in3[34]), .B(inst_cellmath__64_0_in4[34]), .CI(N1710));
ADDFX1 inst_cellmath__64_0_I517 (.CO(N1722), .S(N1721), .A(N1719), .B(N1717), .CI(N1712));
ADDFX1 inst_cellmath__64_0_I518 (.CO(N1724), .S(N1723), .A(inst_cellmath__64_0_in0[47]), .B(N1721), .CI(N1714));
ADDHX1 inst_cellmath__64_0_I519 (.CO(N1726), .S(N1725), .A(inst_cellmath__64_0_in2[35]), .B(inst_cellmath__64_0_in1[35]));
ADDFX1 inst_cellmath__64_0_I520 (.CO(N1728), .S(N1727), .A(inst_cellmath__64_0_in3[35]), .B(inst_cellmath__64_0_in4[35]), .CI(N1718));
ADDFX1 inst_cellmath__64_0_I521 (.CO(N1730), .S(N1729), .A(N1720), .B(N1725), .CI(N1727));
ADDFX1 inst_cellmath__64_0_I522 (.CO(N1732), .S(N1731), .A(N1722), .B(N1729), .CI(inst_cellmath__64_0_in0[48]));
ADDHX1 inst_cellmath__64_0_I523 (.CO(N1734), .S(N1733), .A(inst_cellmath__64_0_in2[36]), .B(inst_cellmath__64_0_in1[36]));
ADDFX1 inst_cellmath__64_0_I524 (.CO(N1736), .S(N1735), .A(inst_cellmath__64_0_in3[36]), .B(inst_cellmath__64_0_in4[36]), .CI(N1726));
ADDFX1 inst_cellmath__64_0_I525 (.CO(N1738), .S(N1737), .A(N1728), .B(N1733), .CI(N1735));
ADDFX1 inst_cellmath__64_0_I526 (.CO(N1740), .S(N1739), .A(N1737), .B(N1730), .CI(inst_cellmath__64_0_in0[49]));
ADDHX1 inst_cellmath__64_0_I527 (.CO(N1742), .S(N1741), .A(inst_cellmath__64_0_in2[37]), .B(inst_cellmath__64_0_in1[37]));
ADDFX1 inst_cellmath__64_0_I528 (.CO(N1744), .S(N1743), .A(inst_cellmath__64_0_in3[37]), .B(inst_cellmath__64_0_in4[37]), .CI(N1734));
ADDFX1 inst_cellmath__64_0_I529 (.CO(N1746), .S(N1745), .A(N1736), .B(N1741), .CI(N1743));
ADDFX1 inst_cellmath__64_0_I530 (.CO(N1748), .S(N1747), .A(N1745), .B(N1738), .CI(inst_cellmath__64_0_in0[50]));
ADDHX1 inst_cellmath__64_0_I531 (.CO(N1750), .S(N1749), .A(inst_cellmath__64_0_in2[38]), .B(inst_cellmath__64_0_in1[38]));
ADDFX1 inst_cellmath__64_0_I532 (.CO(N1752), .S(N1751), .A(inst_cellmath__64_0_in3[38]), .B(inst_cellmath__64_0_in4[38]), .CI(N1742));
ADDFX1 inst_cellmath__64_0_I533 (.CO(N1754), .S(N1753), .A(N1744), .B(N1749), .CI(N1751));
ADDFX1 inst_cellmath__64_0_I534 (.CO(N1756), .S(N1755), .A(N1753), .B(N1746), .CI(inst_cellmath__64_0_in0[51]));
XOR2XL inst_cellmath__64_0_I535 (.Y(N1757), .A(inst_cellmath__64_0_in2[39]), .B(inst_cellmath__64_0_in1[39]));
ADDFX1 inst_cellmath__64_0_I536 (.CO(N1760), .S(N1759), .A(inst_cellmath__64_0_in3[39]), .B(inst_cellmath__64_0_in4[39]), .CI(N1750));
ADDFX1 inst_cellmath__64_0_I537 (.CO(N1762), .S(N1761), .A(N1752), .B(N1757), .CI(N1759));
ADDFX1 inst_cellmath__64_0_I538 (.CO(N1764), .S(N1763), .A(N1761), .B(N1754), .CI(inst_cellmath__64_0_in0[52]));
INVXL inst_cellmath__64_0_I539 (.Y(N1765), .A(N1509));
NOR2XL inst_cellmath__64_0_I540 (.Y(N1767), .A(inst_cellmath__64_0_in3[0]), .B(inst_cellmath__64_0_in2[0]));
NAND2XL inst_cellmath__64_0_I541 (.Y(N1768), .A(inst_cellmath__64_0_in3[0]), .B(inst_cellmath__64_0_in2[0]));
NOR2XL inst_cellmath__64_0_I542 (.Y(N1769), .A(inst_cellmath__64_0_in1[1]), .B(N1513));
NAND2XL inst_cellmath__64_0_I543 (.Y(N1770), .A(inst_cellmath__64_0_in1[1]), .B(N1513));
NOR2XL inst_cellmath__64_0_I544 (.Y(N1771), .A(inst_cellmath__64_0_in1[2]), .B(N1517));
NAND2XL inst_cellmath__64_0_I545 (.Y(N1772), .A(inst_cellmath__64_0_in1[2]), .B(N1517));
NOR2XL inst_cellmath__64_0_I546 (.Y(N1773), .A(inst_cellmath__64_0_in1[3]), .B(N1521));
NAND2XL inst_cellmath__64_0_I547 (.Y(N1774), .A(inst_cellmath__64_0_in1[3]), .B(N1521));
NOR2XL inst_cellmath__64_0_I548 (.Y(N1775), .A(inst_cellmath__64_0_in1[4]), .B(N1525));
NAND2XL inst_cellmath__64_0_I549 (.Y(N1776), .A(inst_cellmath__64_0_in1[4]), .B(N1525));
NOR2XL inst_cellmath__64_0_I550 (.Y(N1777), .A(N1527), .B(N1529));
NAND2XL inst_cellmath__64_0_I551 (.Y(N1778), .A(N1527), .B(N1529));
NOR2XL inst_cellmath__64_0_I552 (.Y(N1779), .A(N1531), .B(N1533));
NAND2XL inst_cellmath__64_0_I553 (.Y(N1780), .A(N1531), .B(N1533));
NOR2XL inst_cellmath__64_0_I554 (.Y(N1781), .A(N1535), .B(N1537));
NAND2XL inst_cellmath__64_0_I555 (.Y(N1782), .A(N1535), .B(N1537));
NOR2X1 inst_cellmath__64_0_I556 (.Y(N1783), .A(N1539), .B(N1541));
NAND2X1 inst_cellmath__64_0_I557 (.Y(N1784), .A(N1539), .B(N1541));
NOR2XL inst_cellmath__64_0_I558 (.Y(N1785), .A(N1542), .B(N1545));
NAND2XL inst_cellmath__64_0_I559 (.Y(N1786), .A(N1542), .B(N1545));
NOR2XL inst_cellmath__64_0_I560 (.Y(N1787), .A(N1546), .B(N1549));
NAND2XL inst_cellmath__64_0_I561 (.Y(N1788), .A(N1546), .B(N1549));
NOR2X1 inst_cellmath__64_0_I562 (.Y(N1789), .A(N1550), .B(N1553));
NAND2X2 inst_cellmath__64_0_I563 (.Y(N1790), .A(N1550), .B(N1553));
NOR2X1 inst_cellmath__64_0_I564 (.Y(N1791), .A(N1554), .B(N1557));
NAND2X2 inst_cellmath__64_0_I565 (.Y(N1792), .A(N1554), .B(N1557));
NOR2XL inst_cellmath__64_0_I566 (.Y(N1793), .A(N1558), .B(N1561));
NAND2XL inst_cellmath__64_0_I567 (.Y(N1794), .A(N1558), .B(N1561));
NOR2XL inst_cellmath__64_0_I568 (.Y(N1795), .A(N1562), .B(N1565));
NAND2XL inst_cellmath__64_0_I569 (.Y(N1796), .A(N1562), .B(N1565));
AOI21XL inst_cellmath__64_0_I572 (.Y(N1799), .A0(N1768), .A1(N1765), .B0(N1767));
INVXL inst_cellmath__64_0_I1430 (.Y(N2875), .A(N1769));
INVXL inst_cellmath__64_0_I1431 (.Y(N2876), .A(N1770));
OAI21XL inst_cellmath__64_0_I580 (.Y(N1807), .A0(N2876), .A1(N1799), .B0(N2875));
AOI21XL inst_cellmath__64_0_I588 (.Y(N1815), .A0(N1772), .A1(N1807), .B0(N1771));
INVXL inst_cellmath__64_0_I1437 (.Y(N2882), .A(N1773));
INVXL inst_cellmath__64_0_I1438 (.Y(N2883), .A(N1774));
OAI21XL inst_cellmath__64_0_I600 (.Y(N1827), .A0(N2883), .A1(N1815), .B0(N2882));
AOI21XL inst_cellmath__64_0_I612 (.Y(N1839), .A0(N1776), .A1(N1827), .B0(N1775));
INVXL inst_cellmath__64_0_I1448 (.Y(N2893), .A(N1777));
INVXL inst_cellmath__64_0_I1449 (.Y(N2894), .A(N1778));
OAI21XL inst_cellmath__64_0_I628 (.Y(N1855), .A0(N2894), .A1(N1839), .B0(N2893));
AOI21XL inst_cellmath__64_0_I644 (.Y(N1871), .A0(N1780), .A1(N1855), .B0(N1779));
INVXL inst_cellmath__64_0_I1463 (.Y(N2908), .A(N1781));
INVXL inst_cellmath__64_0_I1464 (.Y(N2909), .A(N1782));
OAI21XL inst_cellmath__64_0_I664 (.Y(N1891), .A0(N2909), .A1(N1871), .B0(N2908));
AOI21X2 inst_cellmath__64_0_I684 (.Y(N1911), .A0(N1784), .A1(N1891), .B0(N1783));
INVXL inst_cellmath__64_0_I1482 (.Y(N2927), .A(N1785));
INVXL inst_cellmath__64_0_I1483 (.Y(N2928), .A(N1786));
OAI21X2 inst_cellmath__64_0_I708 (.Y(N1935), .A0(N2928), .A1(N1911), .B0(N2927));
AOI21X2 inst_cellmath__64_0_I732 (.Y(N1959), .A0(N1788), .A1(N1935), .B0(N1787));
INVX1 inst_cellmath__64_0_I1505 (.Y(N2950), .A(N1789));
INVX1 inst_cellmath__64_0_I1506 (.Y(N2951), .A(N1790));
OAI21X2 inst_cellmath__64_0_I760 (.Y(N1987), .A0(N2951), .A1(N1959), .B0(N2950));
AOI21X2 inst_cellmath__64_0_I788 (.Y(N2015), .A0(N1792), .A1(N1987), .B0(N1791));
INVXL inst_cellmath__64_0_I1532 (.Y(N2977), .A(N1793));
INVXL inst_cellmath__64_0_I1533 (.Y(N2978), .A(N1794));
OAI21X2 inst_cellmath__64_0_I820 (.Y(N2047), .A0(N2978), .A1(N2015), .B0(N2977));
AOI21X2 inst_cellmath__64_0_I852 (.Y(N2079), .A0(N1796), .A1(N2047), .B0(N1795));
NAND2BXL inst_cellmath__64_0_I875 (.Y(N2102), .AN(N1767), .B(N1768));
NAND2BXL inst_cellmath__64_0_I878 (.Y(N2105), .AN(N1769), .B(N1770));
NAND2BXL inst_cellmath__64_0_I881 (.Y(N2108), .AN(N1771), .B(N1772));
NAND2BXL inst_cellmath__64_0_I884 (.Y(N2111), .AN(N1773), .B(N1774));
NAND2BXL inst_cellmath__64_0_I887 (.Y(N2114), .AN(N1775), .B(N1776));
NAND2BXL inst_cellmath__64_0_I890 (.Y(N2117), .AN(N1777), .B(N1778));
NAND2BXL inst_cellmath__64_0_I893 (.Y(N2120), .AN(N1779), .B(N1780));
NAND2BXL inst_cellmath__64_0_I896 (.Y(N2123), .AN(N1781), .B(N1782));
NAND2BXL inst_cellmath__64_0_I899 (.Y(N2126), .AN(N1783), .B(N1784));
NAND2BXL inst_cellmath__64_0_I902 (.Y(N2129), .AN(N1785), .B(N1786));
NAND2BXL inst_cellmath__64_0_I905 (.Y(N2132), .AN(N1787), .B(N1788));
NAND2BXL inst_cellmath__64_0_I908 (.Y(N2135), .AN(N1789), .B(N1790));
NAND2BXL inst_cellmath__64_0_I911 (.Y(N2138), .AN(N1791), .B(N1792));
NAND2BXL inst_cellmath__64_0_I914 (.Y(N2141), .AN(N1793), .B(N1794));
NAND2BXL inst_cellmath__64_0_I917 (.Y(N2144), .AN(N1795), .B(N1796));
XOR2XL inst_cellmath__64_0_I1669 (.Y(inst_cellmath__64_0_out0[0]), .A(N1765), .B(N2102));
XNOR2X1 inst_cellmath__64_0_I920 (.Y(inst_cellmath__64_0_out0[1]), .A(N1799), .B(N2105));
XOR2XL inst_cellmath__64_0_I1670 (.Y(inst_cellmath__64_0_out0[2]), .A(N1807), .B(N2108));
XNOR2X1 inst_cellmath__64_0_I922 (.Y(inst_cellmath__64_0_out0[3]), .A(N1815), .B(N2111));
XOR2XL inst_cellmath__64_0_I1671 (.Y(inst_cellmath__64_0_out0[4]), .A(N1827), .B(N2114));
XNOR2X1 inst_cellmath__64_0_I924 (.Y(inst_cellmath__64_0_out0[5]), .A(N1839), .B(N2117));
XOR2XL inst_cellmath__64_0_I1672 (.Y(inst_cellmath__64_0_out0[6]), .A(N1855), .B(N2120));
XNOR2X1 inst_cellmath__64_0_I926 (.Y(inst_cellmath__64_0_out0[7]), .A(N1871), .B(N2123));
XOR2XL inst_cellmath__64_0_I1673 (.Y(inst_cellmath__64_0_out0[8]), .A(N1891), .B(N2126));
XNOR2X1 inst_cellmath__64_0_I928 (.Y(inst_cellmath__64_0_out0[9]), .A(N1911), .B(N2129));
XOR2XL inst_cellmath__64_0_I1674 (.Y(inst_cellmath__64_0_out0[10]), .A(N1935), .B(N2132));
XNOR2X1 inst_cellmath__64_0_I930 (.Y(inst_cellmath__64_0_out0[11]), .A(N1959), .B(N2135));
XOR2XL inst_cellmath__64_0_I1675 (.Y(inst_cellmath__64_0_out0[12]), .A(N1987), .B(N2138));
XNOR2X1 inst_cellmath__64_0_I932 (.Y(inst_cellmath__64_0_out0[13]), .A(N2015), .B(N2141));
XOR2XL inst_cellmath__64_0_I1676 (.Y(inst_cellmath__64_0_out0[14]), .A(N2047), .B(N2144));
INVX2 inst_cellmath__64_0_I934 (.Y(N2161), .A(N2079));
NOR2XL inst_cellmath__64_0_I935 (.Y(N2163), .A(N1566), .B(N1571));
NAND2XL inst_cellmath__64_0_I936 (.Y(N2164), .A(N1566), .B(N1571));
NOR2X2 inst_cellmath__64_0_I937 (.Y(N2165), .A(N1572), .B(N1579));
NAND2X1 inst_cellmath__64_0_I938 (.Y(N2166), .A(N1572), .B(N1579));
NOR2X1 inst_cellmath__64_0_I939 (.Y(N2167), .A(N1580), .B(N1587));
NAND2X4 inst_cellmath__64_0_I940 (.Y(N2168), .A(N1580), .B(N1587));
NOR2X1 inst_cellmath__64_0_I941 (.Y(N2169), .A(N1588), .B(N1595));
NAND2X1 inst_cellmath__64_0_I942 (.Y(N2170), .A(N1588), .B(N1595));
NOR2XL inst_cellmath__64_0_I943 (.Y(N2171), .A(N1596), .B(N1603));
NAND2X2 inst_cellmath__64_0_I944 (.Y(N2172), .A(N1596), .B(N1603));
NOR2X1 inst_cellmath__64_0_I945 (.Y(N2173), .A(N1604), .B(N1611));
NAND2X1 inst_cellmath__64_0_I946 (.Y(N2174), .A(N1604), .B(N1611));
NOR2XL inst_cellmath__64_0_I947 (.Y(N2175), .A(N1612), .B(N1619));
NAND2X1 inst_cellmath__64_0_I948 (.Y(N2176), .A(N1612), .B(N1619));
NOR2X1 inst_cellmath__64_0_I949 (.Y(N2177), .A(N1620), .B(N1627));
NAND2X1 inst_cellmath__64_0_I950 (.Y(N2178), .A(N1620), .B(N1627));
NOR2XL inst_cellmath__64_0_I951 (.Y(N2179), .A(N1628), .B(N1635));
NAND2XL inst_cellmath__64_0_I952 (.Y(N2180), .A(N1628), .B(N1635));
NOR2XL inst_cellmath__64_0_I953 (.Y(N2181), .A(N1643), .B(N1636));
NAND2XL inst_cellmath__64_0_I954 (.Y(N2182), .A(N1643), .B(N1636));
NOR2XL inst_cellmath__64_0_I955 (.Y(N2183), .A(N1651), .B(N1644));
NAND2XL inst_cellmath__64_0_I956 (.Y(N2184), .A(N1651), .B(N1644));
NOR2XL inst_cellmath__64_0_I957 (.Y(N2185), .A(N1652), .B(N1659));
NAND2XL inst_cellmath__64_0_I958 (.Y(N2186), .A(N1652), .B(N1659));
NOR2XL inst_cellmath__64_0_I959 (.Y(N2187), .A(N1660), .B(N1667));
NAND2XL inst_cellmath__64_0_I960 (.Y(N2188), .A(N1660), .B(N1667));
NOR2XL inst_cellmath__64_0_I961 (.Y(N2189), .A(N1675), .B(N1668));
NAND2XL inst_cellmath__64_0_I962 (.Y(N2190), .A(N1675), .B(N1668));
NOR2XL inst_cellmath__64_0_I963 (.Y(N2191), .A(N1683), .B(N1676));
NAND2XL inst_cellmath__64_0_I964 (.Y(N2192), .A(N1683), .B(N1676));
NOR2XL inst_cellmath__64_0_I965 (.Y(N2193), .A(N1691), .B(N1684));
NAND2XL inst_cellmath__64_0_I966 (.Y(N2194), .A(N1691), .B(N1684));
NOR2XL inst_cellmath__64_0_I967 (.Y(N2195), .A(N1699), .B(N1692));
NAND2XL inst_cellmath__64_0_I968 (.Y(N2196), .A(N1699), .B(N1692));
NOR2XL inst_cellmath__64_0_I969 (.Y(N2197), .A(N1707), .B(N1700));
NAND2XL inst_cellmath__64_0_I970 (.Y(N2198), .A(N1707), .B(N1700));
NOR2XL inst_cellmath__64_0_I971 (.Y(N2199), .A(N1715), .B(N1708));
NAND2XL inst_cellmath__64_0_I972 (.Y(N2200), .A(N1715), .B(N1708));
NOR2XL inst_cellmath__64_0_I973 (.Y(N2201), .A(N1723), .B(N1716));
NAND2XL inst_cellmath__64_0_I974 (.Y(N2202), .A(N1723), .B(N1716));
NOR2XL inst_cellmath__64_0_I975 (.Y(N2203), .A(N1731), .B(N1724));
NAND2XL inst_cellmath__64_0_I976 (.Y(N2204), .A(N1731), .B(N1724));
NOR2XL inst_cellmath__64_0_I977 (.Y(N2205), .A(N1732), .B(N1739));
NAND2XL inst_cellmath__64_0_I978 (.Y(N2206), .A(N1732), .B(N1739));
NOR2XL inst_cellmath__64_0_I979 (.Y(N2207), .A(N1740), .B(N1747));
NAND2XL inst_cellmath__64_0_I980 (.Y(N2208), .A(N1740), .B(N1747));
NOR2XL inst_cellmath__64_0_I981 (.Y(N2209), .A(N1748), .B(N1755));
NAND2XL inst_cellmath__64_0_I982 (.Y(N2210), .A(N1748), .B(N1755));
AOI21X2 inst_cellmath__64_0_I987 (.Y(N2215), .A0(N2164), .A1(N2161), .B0(N2163));
AOI21X4 inst_cellmath__64_0_I991 (.Y(N2219), .A0(N2168), .A1(N2165), .B0(N2167));
AOI21X1 inst_cellmath__64_0_I995 (.Y(N2223), .A0(N2172), .A1(N2169), .B0(N2171));
AOI21X1 inst_cellmath__64_0_I1003 (.Y(N2231), .A0(N2180), .A1(N2177), .B0(N2179));
AOI21X1 inst_cellmath__64_0_I1007 (.Y(N2235), .A0(N2184), .A1(N2181), .B0(N2183));
NAND2XL inst_cellmath__64_0_I1008 (.Y(N2236), .A(N2184), .B(N2182));
INVXL inst_cellmath__64_0_I1575 (.Y(N3020), .A(N2186));
AOI21XL inst_cellmath__64_0_I1011 (.Y(N2239), .A0(N2188), .A1(N2185), .B0(N2187));
NAND2XL inst_cellmath__64_0_I1012 (.Y(N2240), .A(N2188), .B(N2186));
OAI21XL inst_cellmath__64_0_I1019 (.Y(N2247), .A0(N2240), .A1(N2235), .B0(N2239));
NOR2X1 inst_cellmath__64_0_I1020 (.Y(N2248), .A(N2240), .B(N2236));
AOI21XL inst_cellmath__64_0_I1023 (.Y(N2251), .A0(N2192), .A1(N2189), .B0(N2191));
NAND2XL inst_cellmath__64_0_I1024 (.Y(N2252), .A(N2192), .B(N2190));
INVXL inst_cellmath__64_0_I1583 (.Y(N3028), .A(N2194));
AOI21XL inst_cellmath__64_0_I1027 (.Y(N2255), .A0(N2196), .A1(N2193), .B0(N2195));
NAND2XL inst_cellmath__64_0_I1028 (.Y(N2256), .A(N2196), .B(N2194));
OAI21XL inst_cellmath__64_0_I1035 (.Y(N2263), .A0(N2256), .A1(N2251), .B0(N2255));
NOR2XL inst_cellmath__64_0_I1036 (.Y(N2264), .A(N2256), .B(N2252));
AOI21XL inst_cellmath__64_0_I1039 (.Y(N2267), .A0(N2200), .A1(N2197), .B0(N2199));
NAND2XL inst_cellmath__64_0_I1040 (.Y(N2268), .A(N2200), .B(N2198));
INVXL inst_cellmath__64_0_I1591 (.Y(N3036), .A(N2202));
AOI21XL inst_cellmath__64_0_I1043 (.Y(N2271), .A0(N2204), .A1(N2201), .B0(N2203));
NAND2XL inst_cellmath__64_0_I1044 (.Y(N2272), .A(N2204), .B(N2202));
OAI21XL inst_cellmath__64_0_I1051 (.Y(N2279), .A0(N2272), .A1(N2267), .B0(N2271));
NOR2XL inst_cellmath__64_0_I1052 (.Y(N2280), .A(N2272), .B(N2268));
AOI21XL inst_cellmath__64_0_I1055 (.Y(N2283), .A0(N2208), .A1(N2205), .B0(N2207));
NAND2XL inst_cellmath__64_0_I1056 (.Y(N2284), .A(N2208), .B(N2206));
INVXL inst_cellmath__64_0_I1599 (.Y(N3044), .A(N2210));
INVX2 inst_cellmath__64_0_I1605 (.Y(N3050), .A(N2215));
CLKINVX4 inst_cellmath__64_0_I1608 (.Y(N3053), .A(N2219));
CLKAND2X2 inst_cellmath__64_0_I1680 (.Y(N3054), .A(N2168), .B(N2166));
INVX2 inst_cellmath__64_0_I1612 (.Y(N3057), .A(N2223));
AND2X4 inst_cellmath__64_0_I1682 (.Y(N3060), .A(N2172), .B(N2170));
AO21X1 inst_cellmath__64_0_I2669 (.Y(N3063), .A0(N2176), .A1(N2173), .B0(N2175));
AND2X2 inst_cellmath__64_0_I1684 (.Y(N3066), .A(N2176), .B(N2174));
INVX1 inst_cellmath__64_0_I1624 (.Y(N3069), .A(N2231));
AND2X2 inst_cellmath__64_0_I1686 (.Y(N3072), .A(N2180), .B(N2178));
INVX1 inst_cellmath__64_0_I1628 (.Y(N3073), .A(N3050));
AOI21X4 inst_cellmath__64_0_I1091 (.Y(N2319), .A0(N3054), .A1(N3050), .B0(N3053));
AOI21X4 inst_cellmath__64_0_I1093 (.Y(N2321), .A0(N3060), .A1(N3053), .B0(N3057));
NAND2X4 inst_cellmath__64_0_I1094 (.Y(N2322), .A(N3060), .B(N3054));
AOI21X2 inst_cellmath__64_0_I1095 (.Y(N2323), .A0(N3066), .A1(N3057), .B0(N3063));
NAND2X2 inst_cellmath__64_0_I1096 (.Y(N2324), .A(N3066), .B(N3060));
AOI21X2 inst_cellmath__64_0_I1097 (.Y(N2325), .A0(N3072), .A1(N3063), .B0(N3069));
NAND2X4 inst_cellmath__64_0_I1098 (.Y(N2326), .A(N3072), .B(N3066));
AOI21X2 inst_cellmath__64_0_I1099 (.Y(N2327), .A0(N2248), .A1(N3069), .B0(N2247));
NAND2X2 inst_cellmath__64_0_I1100 (.Y(N2328), .A(N2248), .B(N3072));
AOI21XL inst_cellmath__64_0_I1101 (.Y(N2329), .A0(N2264), .A1(N2247), .B0(N2263));
NAND2X1 inst_cellmath__64_0_I1102 (.Y(N2330), .A(N2264), .B(N2248));
AOI21XL inst_cellmath__64_0_I1103 (.Y(N2331), .A0(N2280), .A1(N2263), .B0(N2279));
NAND2XL inst_cellmath__64_0_I1104 (.Y(N2332), .A(N2280), .B(N2264));
INVXL inst_cellmath__64_0_I1629 (.Y(N3074), .A(N3073));
INVX1 inst_cellmath__64_0_I1630 (.Y(N3075), .A(N2319));
OAI21X4 inst_cellmath__64_0_I1109 (.Y(N2337), .A0(N2322), .A1(N3073), .B0(N2321));
OAI21X4 inst_cellmath__64_0_I1111 (.Y(N2339), .A0(N2324), .A1(N2319), .B0(N2323));
OAI21X2 inst_cellmath__64_0_I1113 (.Y(N2341), .A0(N2326), .A1(N2321), .B0(N2325));
NOR2X2 inst_cellmath__64_0_I1114 (.Y(N2342), .A(N2326), .B(N2322));
OAI21X2 inst_cellmath__64_0_I1115 (.Y(N2343), .A0(N2328), .A1(N2323), .B0(N2327));
NOR2X2 inst_cellmath__64_0_I1116 (.Y(N2344), .A(N2328), .B(N2324));
OAI21X2 inst_cellmath__64_0_I1117 (.Y(N2345), .A0(N2330), .A1(N2325), .B0(N2329));
NOR2X2 inst_cellmath__64_0_I1118 (.Y(N2346), .A(N2330), .B(N2326));
OAI21X1 inst_cellmath__64_0_I1119 (.Y(N2347), .A0(N2332), .A1(N2327), .B0(N2331));
NOR2X2 inst_cellmath__64_0_I1120 (.Y(N2348), .A(N2332), .B(N2328));
INVXL inst_cellmath__64_0_I1631 (.Y(N3076), .A(N3074));
INVXL inst_cellmath__64_0_I1632 (.Y(N3077), .A(N3075));
INVXL inst_cellmath__64_0_I1633 (.Y(N3078), .A(N2337));
INVXL inst_cellmath__64_0_I1634 (.Y(N3079), .A(N2339));
AOI21X2 inst_cellmath__64_0_I1129 (.Y(N2357), .A0(N2342), .A1(N3074), .B0(N2341));
AOI21X2 inst_cellmath__64_0_I1131 (.Y(N2359), .A0(N2344), .A1(N3075), .B0(N2343));
AOI21X4 inst_cellmath__64_0_I1133 (.Y(N2361), .A0(N2346), .A1(N2337), .B0(N2345));
AOI21X4 inst_cellmath__64_0_I1135 (.Y(N2363), .A0(N2348), .A1(N2339), .B0(N2347));
NOR2XL andori2bb1_A_I1756 (.Y(N3114), .A(N3020), .B(N2235));
NOR2XL andori2bb1_A_I1757 (.Y(N3093), .A(N3114), .B(N2185));
NOR2XL andori2bb1_A_I1758 (.Y(N3121), .A(N3028), .B(N2251));
NOR2XL andori2bb1_A_I1759 (.Y(N3099), .A(N3121), .B(N2193));
NOR2XL andori2bb1_A_I1760 (.Y(N3128), .A(N3036), .B(N2267));
NOR2XL andori2bb1_A_I1761 (.Y(N3105), .A(N3128), .B(N2201));
NOR2XL andori2bb1_A_I1762 (.Y(N3135), .A(N3044), .B(N2283));
NOR2XL andori2bb1_A_I1763 (.Y(N3111), .A(N3135), .B(N2209));
NAND2BXL inst_cellmath__64_0_I1204 (.Y(N2432), .AN(N2163), .B(N2164));
NAND2BXL inst_cellmath__64_0_I1207 (.Y(N2435), .AN(N2165), .B(N2166));
NAND2BXL inst_cellmath__64_0_I1210 (.Y(N2438), .AN(N2167), .B(N2168));
NAND2BXL inst_cellmath__64_0_I1213 (.Y(N2441), .AN(N2169), .B(N2170));
NAND2BXL inst_cellmath__64_0_I1216 (.Y(N2444), .AN(N2171), .B(N2172));
NAND2BXL inst_cellmath__64_0_I1219 (.Y(N2447), .AN(N2173), .B(N2174));
NAND2BXL inst_cellmath__64_0_I1222 (.Y(N2450), .AN(N2175), .B(N2176));
NAND2BXL inst_cellmath__64_0_I1225 (.Y(N2453), .AN(N2177), .B(N2178));
NAND2BXL inst_cellmath__64_0_I1228 (.Y(N2456), .AN(N2179), .B(N2180));
NAND2BXL inst_cellmath__64_0_I1231 (.Y(N2459), .AN(N2181), .B(N2182));
NAND2BXL inst_cellmath__64_0_I1234 (.Y(N2462), .AN(N2183), .B(N2184));
NAND2BXL inst_cellmath__64_0_I1237 (.Y(N2680), .AN(N2185), .B(N2186));
NAND2BXL inst_cellmath__64_0_I1240 (.Y(N2691), .AN(N2187), .B(N2188));
NAND2BXL inst_cellmath__64_0_I1243 (.Y(N2471), .AN(N2189), .B(N2190));
NAND2BXL inst_cellmath__64_0_I1246 (.Y(N2474), .AN(N2191), .B(N2192));
NAND2BXL inst_cellmath__64_0_I1249 (.Y(N2709), .AN(N2193), .B(N2194));
NAND2BXL inst_cellmath__64_0_I1252 (.Y(N2720), .AN(N2195), .B(N2196));
NAND2BXL inst_cellmath__64_0_I1255 (.Y(N2483), .AN(N2197), .B(N2198));
NAND2BXL inst_cellmath__64_0_I1258 (.Y(N2486), .AN(N2199), .B(N2200));
NAND2BXL inst_cellmath__64_0_I1261 (.Y(N2738), .AN(N2201), .B(N2202));
NAND2BXL inst_cellmath__64_0_I1264 (.Y(N2749), .AN(N2203), .B(N2204));
NAND2BXL inst_cellmath__64_0_I1267 (.Y(N2495), .AN(N2205), .B(N2206));
NAND2BXL inst_cellmath__64_0_I1270 (.Y(N2498), .AN(N2207), .B(N2208));
NAND2BXL inst_cellmath__64_0_I1273 (.Y(N2767), .AN(N2209), .B(N2210));
XNOR2X1 inst_cellmath__64_0_I1731 (.Y(N2778), .A(N1763), .B(N1756));
XOR2XL inst_cellmath__64_0_I1696 (.Y(inst_cellmath__64_0_out0[15]), .A(N2161), .B(N2432));
XNOR2X1 inst_cellmath__64_0_I1279 (.Y(inst_cellmath__64_0_out0[16]), .A(N3076), .B(N2435));
XNOR2X1 inst_cellmath__64_0_I1280 (.Y(inst_cellmath__64_0_out0[18]), .A(N3077), .B(N2441));
XNOR2X1 inst_cellmath__64_0_I2670 (.Y(inst_cellmath__64_0_out0[20]), .A(N3078), .B(N2447));
XNOR2X1 inst_cellmath__64_0_I2671 (.Y(inst_cellmath__64_0_out0[22]), .A(N3079), .B(N2453));
XNOR2X1 inst_cellmath__64_0_I2672 (.Y(inst_cellmath__64_0_out0[24]), .A(N2357), .B(N2459));
XNOR2XL inst_cellmath__64_0_I2673 (.Y(inst_cellmath__64_0_out0[28]), .A(N2359), .B(N2471));
XNOR2X1 inst_cellmath__64_0_I2674 (.Y(inst_cellmath__64_0_out0[32]), .A(N2361), .B(N2483));
XNOR2X1 inst_cellmath__64_0_I2675 (.Y(inst_cellmath__64_0_out0[36]), .A(N2495), .B(N2363));
XOR2XL node_cs_reduced_ii_local_A_I1701 (.Y(N2516), .A(N2438), .B(N2166));
XOR2XL node_cs_reduced_ii_local_A_I1702 (.Y(N2515), .A(N2438), .B(N2165));
MX2XL inst_cellmath__64_0_I1288 (.Y(inst_cellmath__64_0_out0[17]), .A(N2516), .B(N2515), .S0(N3076));
XOR2XL node_cs_reduced_ii_local_A_I1703 (.Y(N2519), .A(N2170), .B(N2444));
XOR2XL node_cs_reduced_ii_local_A_I1704 (.Y(N2518), .A(N2444), .B(N2169));
MX2XL inst_cellmath__64_0_I1290 (.Y(inst_cellmath__64_0_out0[19]), .A(N2519), .B(N2518), .S0(N3077));
XOR2XL node_cs_reduced_ii_local_A_I1705 (.Y(N2522), .A(N2174), .B(N2450));
XOR2XL node_cs_reduced_ii_local_A_I1706 (.Y(N2521), .A(N2450), .B(N2173));
MX2XL inst_cellmath__64_0_I1292 (.Y(inst_cellmath__64_0_out0[21]), .A(N2522), .B(N2521), .S0(N3078));
XOR2XL node_cs_reduced_ii_local_A_I1707 (.Y(N2525), .A(N2456), .B(N2178));
XOR2XL node_cs_reduced_ii_local_A_I1708 (.Y(N2524), .A(N2456), .B(N2177));
MX2XL inst_cellmath__64_0_I1294 (.Y(inst_cellmath__64_0_out0[23]), .A(N2525), .B(N2524), .S0(N3079));
XOR2XL node_cs_reduced_ii_local_A_I1709 (.Y(N2528), .A(N2462), .B(N2182));
XOR2XL node_cs_reduced_ii_local_A_I1710 (.Y(N2527), .A(N2462), .B(N2181));
MX2XL inst_cellmath__64_0_I1296 (.Y(inst_cellmath__64_0_out0[25]), .A(N2528), .B(N2527), .S0(N2357));
XOR2XL node_cs_ii_local_alt_A_I1362 (.Y(N2530), .A(N2680), .B(N2235));
NAND2XL node_cs_ii_local_alt_A_I1363 (.Y(N2678), .A(N2236), .B(N2235));
XNOR2X1 node_cs_ii_local_alt_A_I1364 (.Y(N2531), .A(N2680), .B(N2678));
MXI2XL inst_cellmath__64_0_I1298 (.Y(inst_cellmath__64_0_out0[26]), .A(N2531), .B(N2530), .S0(N2357));
XOR2XL node_cs_ii_local_alt_A_I1366 (.Y(N2533), .A(N2691), .B(N3093));
OAI21XL node_cs_ii_local_alt_A_I1711 (.Y(N2689), .A0(N3020), .A1(N2236), .B0(N3093));
XNOR2X1 node_cs_ii_local_alt_A_I1368 (.Y(N2534), .A(N2691), .B(N2689));
MXI2XL inst_cellmath__64_0_I1300 (.Y(inst_cellmath__64_0_out0[27]), .A(N2534), .B(N2533), .S0(N2357));
XOR2XL node_cs_reduced_ii_local_A_I1712 (.Y(N2537), .A(N2474), .B(N2190));
XOR2XL node_cs_reduced_ii_local_A_I1713 (.Y(N2536), .A(N2474), .B(N2189));
MX2XL inst_cellmath__64_0_I2676 (.Y(inst_cellmath__64_0_out0[29]), .A(N2537), .B(N2536), .S0(N2359));
XOR2XL node_cs_ii_local_alt_A_I1372 (.Y(N2539), .A(N2709), .B(N2251));
NAND2XL node_cs_ii_local_alt_A_I1373 (.Y(N2707), .A(N2252), .B(N2251));
XNOR2X1 node_cs_ii_local_alt_A_I1374 (.Y(N2540), .A(N2709), .B(N2707));
MXI2XL inst_cellmath__64_0_I1304 (.Y(inst_cellmath__64_0_out0[30]), .A(N2540), .B(N2539), .S0(N2359));
XOR2XL node_cs_ii_local_alt_A_I1376 (.Y(N2542), .A(N2720), .B(N3099));
OAI21XL node_cs_ii_local_alt_A_I1714 (.Y(N2718), .A0(N3028), .A1(N2252), .B0(N3099));
XNOR2X1 node_cs_ii_local_alt_A_I1378 (.Y(N2543), .A(N2720), .B(N2718));
MXI2XL inst_cellmath__64_0_I1306 (.Y(inst_cellmath__64_0_out0[31]), .A(N2543), .B(N2542), .S0(N2359));
XOR2XL node_cs_reduced_ii_local_A_I1715 (.Y(N2546), .A(N2486), .B(N2198));
XOR2XL node_cs_reduced_ii_local_A_I1716 (.Y(N2545), .A(N2486), .B(N2197));
MX2XL inst_cellmath__64_0_I2677 (.Y(inst_cellmath__64_0_out0[33]), .A(N2546), .B(N2545), .S0(N2361));
XOR2XL node_cs_ii_local_alt_A_I1382 (.Y(N2548), .A(N2738), .B(N2267));
NAND2XL node_cs_ii_local_alt_A_I1383 (.Y(N2736), .A(N2268), .B(N2267));
XNOR2X1 node_cs_ii_local_alt_A_I1384 (.Y(N2549), .A(N2738), .B(N2736));
MXI2XL inst_cellmath__64_0_I1310 (.Y(inst_cellmath__64_0_out0[34]), .A(N2549), .B(N2548), .S0(N2361));
XOR2XL node_cs_ii_local_alt_A_I1386 (.Y(N2551), .A(N2749), .B(N3105));
OAI21XL node_cs_ii_local_alt_A_I1717 (.Y(N2747), .A0(N3036), .A1(N2268), .B0(N3105));
XNOR2X1 node_cs_ii_local_alt_A_I1388 (.Y(N2552), .A(N2749), .B(N2747));
MXI2XL inst_cellmath__64_0_I1312 (.Y(inst_cellmath__64_0_out0[35]), .A(N2552), .B(N2551), .S0(N2361));
XOR2XL node_cs_reduced_ii_local_A_I1718 (.Y(N2555), .A(N2498), .B(N2206));
XOR2XL node_cs_reduced_ii_local_A_I1719 (.Y(N2554), .A(N2498), .B(N2205));
MX2XL inst_cellmath__64_0_I1314 (.Y(inst_cellmath__64_0_out0[37]), .A(N2555), .B(N2554), .S0(N2363));
XOR2XL node_cs_ii_local_alt_A_I1392 (.Y(N2557), .A(N2767), .B(N2283));
NAND2XL node_cs_ii_local_alt_A_I1393 (.Y(N2765), .A(N2284), .B(N2283));
XNOR2X1 node_cs_ii_local_alt_A_I1394 (.Y(N2558), .A(N2767), .B(N2765));
MXI2XL inst_cellmath__64_0_I1316 (.Y(inst_cellmath__64_0_out0[38]), .A(N2558), .B(N2557), .S0(N2363));
XOR2XL node_cs_ii_local_alt_A_I1396 (.Y(N2560), .A(N2778), .B(N3111));
OAI21XL node_cs_ii_local_alt_A_I1720 (.Y(N2776), .A0(N3044), .A1(N2284), .B0(N3111));
XNOR2X1 node_cs_ii_local_alt_A_I1398 (.Y(N2561), .A(N2778), .B(N2776));
MXI2XL inst_cellmath__64_0_I1318 (.Y(inst_cellmath__64_0_out0[39]), .A(N2561), .B(N2560), .S0(N2363));
endmodule

module cynw_cm_float_rcp_inst_cellmath__68_0_bdw1471647203_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1,
	inst_cellmath__68_0_in2
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__68_0_out0;
input  inst_cellmath__68_0_in0;
input [39:17] inst_cellmath__68_0_in1;
input  inst_cellmath__68_0_in2;
wire N50,N51,N52,N53,N54,N55,N56 
	,N57,N58,N59,N60,N61,N62,N63,N64 
	,N65,N66,N67,N68,N69,N70,N71,N72 
	,N122,N137;
INVXL inst_cellmath__68_0_I0 (.Y(N50), .A(inst_cellmath__68_0_in1[17]));
INVXL inst_cellmath__68_0_I1 (.Y(N51), .A(inst_cellmath__68_0_in1[18]));
INVXL inst_cellmath__68_0_I2 (.Y(N52), .A(inst_cellmath__68_0_in1[19]));
INVXL inst_cellmath__68_0_I3 (.Y(N53), .A(inst_cellmath__68_0_in1[20]));
INVXL inst_cellmath__68_0_I4 (.Y(N54), .A(inst_cellmath__68_0_in1[21]));
INVXL inst_cellmath__68_0_I5 (.Y(N55), .A(inst_cellmath__68_0_in1[22]));
INVXL inst_cellmath__68_0_I6 (.Y(N56), .A(inst_cellmath__68_0_in1[23]));
INVXL inst_cellmath__68_0_I7 (.Y(N57), .A(inst_cellmath__68_0_in1[24]));
INVXL inst_cellmath__68_0_I8 (.Y(N58), .A(inst_cellmath__68_0_in1[25]));
INVXL inst_cellmath__68_0_I9 (.Y(N59), .A(inst_cellmath__68_0_in1[26]));
INVXL inst_cellmath__68_0_I10 (.Y(N60), .A(inst_cellmath__68_0_in1[27]));
INVXL inst_cellmath__68_0_I11 (.Y(N61), .A(inst_cellmath__68_0_in1[28]));
INVXL inst_cellmath__68_0_I12 (.Y(N62), .A(inst_cellmath__68_0_in1[29]));
INVXL inst_cellmath__68_0_I13 (.Y(N63), .A(inst_cellmath__68_0_in1[30]));
INVXL inst_cellmath__68_0_I14 (.Y(N64), .A(inst_cellmath__68_0_in1[31]));
INVXL inst_cellmath__68_0_I15 (.Y(N65), .A(inst_cellmath__68_0_in1[32]));
INVXL inst_cellmath__68_0_I16 (.Y(N66), .A(inst_cellmath__68_0_in1[33]));
INVXL inst_cellmath__68_0_I17 (.Y(N67), .A(inst_cellmath__68_0_in1[34]));
INVXL inst_cellmath__68_0_I18 (.Y(N68), .A(inst_cellmath__68_0_in1[35]));
INVXL inst_cellmath__68_0_I19 (.Y(N69), .A(inst_cellmath__68_0_in1[36]));
INVXL inst_cellmath__68_0_I20 (.Y(N70), .A(inst_cellmath__68_0_in1[37]));
INVXL inst_cellmath__68_0_I21 (.Y(N71), .A(inst_cellmath__68_0_in1[38]));
INVXL inst_cellmath__68_0_I22 (.Y(N72), .A(inst_cellmath__68_0_in1[39]));
INVXL inst_cellmath__68_0_I71 (.Y(N122), .A(inst_cellmath__68_0_in2));
INVXL inst_cellmath__68_0_I86 (.Y(N137), .A(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I47 (.Y(inst_cellmath__68_0_out0[0]), .A0(N137), .A1(N122), .B0(N50), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I48 (.Y(inst_cellmath__68_0_out0[1]), .A0(N137), .A1(N122), .B0(N51), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I49 (.Y(inst_cellmath__68_0_out0[2]), .A0(N137), .A1(N122), .B0(N52), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I50 (.Y(inst_cellmath__68_0_out0[3]), .A0(N137), .A1(N122), .B0(N53), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I51 (.Y(inst_cellmath__68_0_out0[4]), .A0(N137), .A1(N122), .B0(N54), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I52 (.Y(inst_cellmath__68_0_out0[5]), .A0(N137), .A1(N122), .B0(N55), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I53 (.Y(inst_cellmath__68_0_out0[6]), .A0(N137), .A1(N122), .B0(N56), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I54 (.Y(inst_cellmath__68_0_out0[7]), .A0(N137), .A1(N122), .B0(N57), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I55 (.Y(inst_cellmath__68_0_out0[8]), .A0(N137), .A1(N122), .B0(N58), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I56 (.Y(inst_cellmath__68_0_out0[9]), .A0(N137), .A1(N122), .B0(N59), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I57 (.Y(inst_cellmath__68_0_out0[10]), .A0(N137), .A1(N122), .B0(N60), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I58 (.Y(inst_cellmath__68_0_out0[11]), .A0(N137), .A1(N122), .B0(N61), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I59 (.Y(inst_cellmath__68_0_out0[12]), .A0(N137), .A1(N122), .B0(N62), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I60 (.Y(inst_cellmath__68_0_out0[13]), .A0(N137), .A1(N122), .B0(N63), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I61 (.Y(inst_cellmath__68_0_out0[14]), .A0(N137), .A1(N122), .B0(N64), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I62 (.Y(inst_cellmath__68_0_out0[15]), .A0(N137), .A1(N122), .B0(N65), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I63 (.Y(inst_cellmath__68_0_out0[16]), .A0(N122), .A1(N137), .B0(N66), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I64 (.Y(inst_cellmath__68_0_out0[17]), .A0(N137), .A1(N122), .B0(N67), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I65 (.Y(inst_cellmath__68_0_out0[18]), .A0(N137), .A1(N122), .B0(N68), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I66 (.Y(inst_cellmath__68_0_out0[19]), .A0(N137), .A1(N122), .B0(N69), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I67 (.Y(inst_cellmath__68_0_out0[20]), .A0(N137), .A1(N122), .B0(N70), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I68 (.Y(inst_cellmath__68_0_out0[21]), .A0(N137), .A1(N122), .B0(N71), .B1(inst_cellmath__68_0_in0));
AOI22XL inst_cellmath__68_0_I69 (.Y(inst_cellmath__68_0_out0[22]), .A0(N137), .A1(N122), .B0(N72), .B1(inst_cellmath__68_0_in0));
endmodule

/* CADENCE  uLb2TQrfqho= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



