/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:28 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417;
wire N4032,N8724,N8762,N8769,N8776,N8782,N8785 
	,N8794,N8803,N8812,N8821,N8830,N8839,N8848,N8857 
	,N8866,N8875,N8884,N8893,N8902,N8911,N8920,N8929 
	,N8938,N8947,N8956,N8965,N9174,N9179,N9184,N9189 
	,N9194,N9199,N9204,N9209,N9214,N9219,N9224,N9229 
	,N9234,N9239,N9244,N9249,N9254,N9259,N9264,N9269 
	,N9274,N9279,N9467,N9505,N9507,N9512,N9514,N9540 
	,N9566,N9592,N9759,N9765,N9768,N9777,N9786,N9795 
	,N9804,N9813,N9822,N9831,N9840,N9849,N9858,N9867 
	,N9876,N9885,N9894,N9903,N9912,N9921,N9930,N9939 
	,N9948,N9957,N9963,N9966,N9972,N9975,N9981,N9984 
	,N9990,N9993,N9999,N10002,N10008,N10011,N10017,N10020 
	,N10026,N10029,N10035,N10038,N10044,N10047,N10053,N10056 
	,N10062,N10065,N10071,N10074,N10080,N10083,N10089,N10092 
	,N10098,N10101,N10107,N10110,N10116,N10119,N10125,N10128 
	,N10134,N10137,N10143,N10146,N10152,N10157,N10162,N10167 
	,N10172,N10177,N10182,N10187,N10192,N10197,N10202,N10207 
	,N10212,N10217,N10222,N10227,N10232,N10237,N10242,N10247 
	,N10252,N10257,N10262,N10412,N10438,N10464,N10490,N10581 
	,N10583,N10616,N10621,N10623,N10625,N10627,N10630,N10632 
	,N10637,N10639,N10643,N10694,N10696,N10703,N10705,N10712 
	,N10714,N10721,N10723,N10730,N10732,N10739,N10741,N10748 
	,N10750,N10757,N10759,N10766,N10768,N10774,N10776,N10827 
	,N10829,N10831,N10845,N10847,N10872,N11135,N11141,N11147 
	,N11153,N11159,N11165,N11171,N11177,N11239,N11241,N11343 
	,N11345,N11350,N11352,N11357,N11359,N11364,N11366,N11373 
	,N11378,N11385,N11387,N11392,N11401,N11406,N11408,N11425 
	,N11432,N11447,N11449,N11454,N11468,N11470,N11475,N11500 
	,N11506,N11512,N11518,N11524,N11530,N11536,N11542,N11548 
	,N11554,N11560,N11564,N11566,N11570,N11572,N11675,N11678 
	,N11686,N11694,N11702,N11710,N11718,N11726,N11734,N11742 
	,N11750,N11758,N11766,N11774,N11782,N11790,N11798,N11806 
	,N11814,N11822,N11830,N12999,N13000,N13001,N13002,N13003 
	,N13004;
reg x_reg_L0_21__retimed_I6170_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6170_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908;
	end
assign N11830 = x_reg_L0_21__retimed_I6170_QOUT;
reg x_reg_L0_21__retimed_I6167_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6167_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168;
	end
assign N11822 = x_reg_L0_21__retimed_I6167_QOUT;
reg x_reg_L0_21__retimed_I6164_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6164_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985;
	end
assign N11814 = x_reg_L0_21__retimed_I6164_QOUT;
reg x_reg_L0_21__retimed_I6161_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6161_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250;
	end
assign N11806 = x_reg_L0_21__retimed_I6161_QOUT;
reg x_reg_L0_21__retimed_I6158_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6158_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069;
	end
assign N11798 = x_reg_L0_21__retimed_I6158_QOUT;
reg x_reg_L0_21__retimed_I6155_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6155_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336;
	end
assign N11790 = x_reg_L0_21__retimed_I6155_QOUT;
reg x_reg_L0_21__retimed_I6152_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6152_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154;
	end
assign N11782 = x_reg_L0_21__retimed_I6152_QOUT;
reg x_reg_L0_21__retimed_I6149_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6149_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413;
	end
assign N11774 = x_reg_L0_21__retimed_I6149_QOUT;
reg x_reg_L0_21__retimed_I6146_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6146_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233;
	end
assign N11766 = x_reg_L0_21__retimed_I6146_QOUT;
reg x_reg_L0_21__retimed_I6143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6143_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501;
	end
assign N11758 = x_reg_L0_21__retimed_I6143_QOUT;
reg x_reg_L0_21__retimed_I6140_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6140_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320;
	end
assign N11750 = x_reg_L0_21__retimed_I6140_QOUT;
reg x_reg_L0_21__retimed_I6137_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6137_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591;
	end
assign N11742 = x_reg_L0_21__retimed_I6137_QOUT;
reg x_reg_L0_21__retimed_I6134_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6134_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407;
	end
assign N11734 = x_reg_L0_21__retimed_I6134_QOUT;
reg x_reg_L0_21__retimed_I6131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6131_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672;
	end
assign N11726 = x_reg_L0_21__retimed_I6131_QOUT;
reg x_reg_L0_21__retimed_I6128_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6128_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475;
	end
assign N11718 = x_reg_L0_21__retimed_I6128_QOUT;
reg x_reg_L0_21__retimed_I6125_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6125_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755;
	end
assign N11710 = x_reg_L0_21__retimed_I6125_QOUT;
reg x_reg_L0_21__retimed_I6122_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6122_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561;
	end
assign N11702 = x_reg_L0_21__retimed_I6122_QOUT;
reg x_reg_L0_21__retimed_I6119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6119_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840;
	end
assign N11694 = x_reg_L0_21__retimed_I6119_QOUT;
reg x_reg_L0_21__retimed_I6116_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6116_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645;
	end
assign N11686 = x_reg_L0_21__retimed_I6116_QOUT;
reg x_reg_L0_21__retimed_I6113_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6113_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917;
	end
assign N11678 = x_reg_L0_21__retimed_I6113_QOUT;
reg x_reg_L0_21__retimed_I6112_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6112_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178;
	end
assign N11675 = x_reg_L0_21__retimed_I6112_QOUT;
reg x_reg_L0_21__retimed_I6090_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6090_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934;
	end
assign N11572 = x_reg_L0_21__retimed_I6090_QOUT;
reg x_reg_L0_21__retimed_I6089_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6089_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254;
	end
assign N11570 = x_reg_L0_21__retimed_I6089_QOUT;
reg x_reg_L0_21__retimed_I6088_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6088_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604;
	end
assign N11566 = x_reg_L0_21__retimed_I6088_QOUT;
reg x_reg_L0_21__retimed_I6087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6087_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144;
	end
assign N11564 = x_reg_L0_21__retimed_I6087_QOUT;
reg x_reg_L0_21__retimed_I6086_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6086_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734;
	end
assign N11560 = x_reg_L0_21__retimed_I6086_QOUT;
reg x_reg_L0_21__retimed_I6084_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6084_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414;
	end
assign N11554 = x_reg_L0_21__retimed_I6084_QOUT;
reg x_reg_L0_21__retimed_I6082_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6082_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538;
	end
assign N11548 = x_reg_L0_21__retimed_I6082_QOUT;
reg x_reg_L0_21__retimed_I6080_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6080_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209;
	end
assign N11542 = x_reg_L0_21__retimed_I6080_QOUT;
reg x_reg_L0_21__retimed_I6078_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6078_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339;
	end
assign N11536 = x_reg_L0_21__retimed_I6078_QOUT;
reg x_reg_L0_21__retimed_I6076_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6076_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014;
	end
assign N11530 = x_reg_L0_21__retimed_I6076_QOUT;
reg x_reg_L0_21__retimed_I6074_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6074_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682;
	end
assign N11524 = x_reg_L0_21__retimed_I6074_QOUT;
reg x_reg_L0_21__retimed_I6072_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6072_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821;
	end
assign N11518 = x_reg_L0_21__retimed_I6072_QOUT;
reg x_reg_L0_21__retimed_I6070_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6070_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483;
	end
assign N11512 = x_reg_L0_21__retimed_I6070_QOUT;
reg x_reg_L0_21__retimed_I6068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6068_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617;
	end
assign N11506 = x_reg_L0_21__retimed_I6068_QOUT;
reg x_reg_L0_21__retimed_I6066_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6066_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293;
	end
assign N11500 = x_reg_L0_21__retimed_I6066_QOUT;
reg x_reg_L0_21__retimed_I6056_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6056_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0];
	end
assign N11475 = x_reg_L0_21__retimed_I6056_QOUT;
reg x_reg_L0_21__retimed_I6054_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6054_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18];
	end
assign N11470 = x_reg_L0_21__retimed_I6054_QOUT;
reg x_reg_L0_21__retimed_I6053_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6053_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17];
	end
assign N11468 = x_reg_L0_21__retimed_I6053_QOUT;
reg x_reg_L0_21__retimed_I6047_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6047_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19];
	end
assign N11454 = x_reg_L0_21__retimed_I6047_QOUT;
reg x_reg_L0_21__retimed_I6045_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6045_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21];
	end
assign N11449 = x_reg_L0_21__retimed_I6045_QOUT;
reg x_reg_L0_21__retimed_I6044_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6044_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20];
	end
assign N11447 = x_reg_L0_21__retimed_I6044_QOUT;
reg x_reg_L1_21__retimed_I6038_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6038_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1];
	end
assign N11432 = x_reg_L1_21__retimed_I6038_QOUT;
reg x_reg_L1_21__retimed_I6035_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I6035_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6];
	end
assign N11425 = x_reg_L1_21__retimed_I6035_QOUT;
reg x_reg_L0_21__retimed_I6028_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6028_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12];
	end
assign N11408 = x_reg_L0_21__retimed_I6028_QOUT;
reg x_reg_L0_21__retimed_I6027_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6027_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11];
	end
assign N11406 = x_reg_L0_21__retimed_I6027_QOUT;
reg x_reg_L0_21__retimed_I6025_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6025_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7];
	end
assign N11401 = x_reg_L0_21__retimed_I6025_QOUT;
reg x_reg_L0_21__retimed_I6021_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6021_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3];
	end
assign N11392 = x_reg_L0_21__retimed_I6021_QOUT;
reg x_reg_L0_21__retimed_I6019_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6019_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14];
	end
assign N11387 = x_reg_L0_21__retimed_I6019_QOUT;
reg x_reg_L0_21__retimed_I6018_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6018_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13];
	end
assign N11385 = x_reg_L0_21__retimed_I6018_QOUT;
reg x_reg_L0_21__retimed_I6015_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6015_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8];
	end
assign N11378 = x_reg_L0_21__retimed_I6015_QOUT;
reg x_reg_L0_21__retimed_I6013_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6013_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6];
	end
assign N11373 = x_reg_L0_21__retimed_I6013_QOUT;
reg x_reg_L0_21__retimed_I6010_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6010_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10];
	end
assign N11366 = x_reg_L0_21__retimed_I6010_QOUT;
reg x_reg_L0_21__retimed_I6009_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6009_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9];
	end
assign N11364 = x_reg_L0_21__retimed_I6009_QOUT;
reg x_reg_L0_21__retimed_I6007_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6007_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5];
	end
assign N11359 = x_reg_L0_21__retimed_I6007_QOUT;
reg x_reg_L0_21__retimed_I6006_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6006_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4];
	end
assign N11357 = x_reg_L0_21__retimed_I6006_QOUT;
reg x_reg_L0_21__retimed_I6004_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6004_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2];
	end
assign N11352 = x_reg_L0_21__retimed_I6004_QOUT;
reg x_reg_L0_21__retimed_I6003_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6003_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1];
	end
assign N11350 = x_reg_L0_21__retimed_I6003_QOUT;
reg x_reg_L0_21__retimed_I6001_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6001_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16];
	end
assign N11345 = x_reg_L0_21__retimed_I6001_QOUT;
reg x_reg_L0_21__retimed_I6000_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I6000_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15];
	end
assign N11343 = x_reg_L0_21__retimed_I6000_QOUT;
reg x_reg_L0_21__retimed_I5966_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5966_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25];
	end
assign N11241 = x_reg_L0_21__retimed_I5966_QOUT;
reg x_reg_L0_21__retimed_I5965_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5965_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24];
	end
assign N11239 = x_reg_L0_21__retimed_I5965_QOUT;
reg x_reg_L0_21__retimed_I5945_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5945_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415;
	end
assign N11177 = x_reg_L0_21__retimed_I5945_QOUT;
reg x_reg_L0_21__retimed_I5943_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5943_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100;
	end
assign N11171 = x_reg_L0_21__retimed_I5943_QOUT;
reg x_reg_L0_21__retimed_I5941_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5941_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219;
	end
assign N11165 = x_reg_L0_21__retimed_I5941_QOUT;
reg x_reg_L0_21__retimed_I5939_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5939_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900;
	end
assign N11159 = x_reg_L0_21__retimed_I5939_QOUT;
reg x_reg_L0_21__retimed_I5937_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5937_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571;
	end
assign N11153 = x_reg_L0_21__retimed_I5937_QOUT;
reg x_reg_L0_21__retimed_I5935_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5935_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704;
	end
assign N11147 = x_reg_L0_21__retimed_I5935_QOUT;
reg x_reg_L0_21__retimed_I5933_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5933_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379;
	end
assign N11141 = x_reg_L0_21__retimed_I5933_QOUT;
reg x_reg_L0_21__retimed_I5931_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5931_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503;
	end
assign N11135 = x_reg_L0_21__retimed_I5931_QOUT;
reg x_reg_L0_21__retimed_I5845_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5845_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4;
	end
assign N10872 = x_reg_L0_21__retimed_I5845_QOUT;
reg x_reg_L0_21__retimed_I5838_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5838_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23];
	end
assign N10847 = x_reg_L0_21__retimed_I5838_QOUT;
reg x_reg_L0_21__retimed_I5837_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5837_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22];
	end
assign N10845 = x_reg_L0_21__retimed_I5837_QOUT;
reg x_reg_L0_21__retimed_I5831_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5831_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446;
	end
assign N10831 = x_reg_L0_21__retimed_I5831_QOUT;
reg x_reg_L0_21__retimed_I5830_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5830_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445;
	end
assign N10829 = x_reg_L0_21__retimed_I5830_QOUT;
reg x_reg_L0_21__retimed_I5829_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5829_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8;
	end
assign N10827 = x_reg_L0_21__retimed_I5829_QOUT;
reg x_reg_L0_21__retimed_I5813_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5813_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8];
	end
assign N10776 = x_reg_L0_21__retimed_I5813_QOUT;
reg x_reg_L0_21__retimed_I5812_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5812_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8];
	end
assign N10774 = x_reg_L0_21__retimed_I5812_QOUT;
reg x_reg_L0_21__retimed_I5810_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5810_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1];
	end
assign N10768 = x_reg_L0_21__retimed_I5810_QOUT;
reg x_reg_L0_21__retimed_I5809_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5809_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1];
	end
assign N10766 = x_reg_L0_21__retimed_I5809_QOUT;
reg x_reg_L0_21__retimed_I5807_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5807_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3];
	end
assign N10759 = x_reg_L0_21__retimed_I5807_QOUT;
reg x_reg_L0_21__retimed_I5806_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5806_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3];
	end
assign N10757 = x_reg_L0_21__retimed_I5806_QOUT;
reg x_reg_L0_21__retimed_I5804_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5804_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6];
	end
assign N10750 = x_reg_L0_21__retimed_I5804_QOUT;
reg x_reg_L0_21__retimed_I5803_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5803_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6];
	end
assign N10748 = x_reg_L0_21__retimed_I5803_QOUT;
reg x_reg_L0_21__retimed_I5801_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5801_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
	end
assign N10741 = x_reg_L0_21__retimed_I5801_QOUT;
reg x_reg_L0_21__retimed_I5800_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5800_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7];
	end
assign N10739 = x_reg_L0_21__retimed_I5800_QOUT;
reg x_reg_L0_21__retimed_I5798_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5798_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9];
	end
assign N10732 = x_reg_L0_21__retimed_I5798_QOUT;
reg x_reg_L0_21__retimed_I5797_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5797_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9];
	end
assign N10730 = x_reg_L0_21__retimed_I5797_QOUT;
reg x_reg_L0_21__retimed_I5795_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5795_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5];
	end
assign N10723 = x_reg_L0_21__retimed_I5795_QOUT;
reg x_reg_L0_21__retimed_I5794_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5794_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5];
	end
assign N10721 = x_reg_L0_21__retimed_I5794_QOUT;
reg x_reg_L0_21__retimed_I5792_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5792_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4];
	end
assign N10714 = x_reg_L0_21__retimed_I5792_QOUT;
reg x_reg_L0_21__retimed_I5791_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5791_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4];
	end
assign N10712 = x_reg_L0_21__retimed_I5791_QOUT;
reg x_reg_L0_21__retimed_I5789_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5789_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2];
	end
assign N10705 = x_reg_L0_21__retimed_I5789_QOUT;
reg x_reg_L0_21__retimed_I5788_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5788_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2];
	end
assign N10703 = x_reg_L0_21__retimed_I5788_QOUT;
reg x_reg_L0_21__retimed_I5786_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5786_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0];
	end
assign N10696 = x_reg_L0_21__retimed_I5786_QOUT;
reg x_reg_L0_21__retimed_I5785_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5785_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0];
	end
assign N10694 = x_reg_L0_21__retimed_I5785_QOUT;
reg x_reg_L1_21__retimed_I5765_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5765_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9];
	end
assign N10643 = x_reg_L1_21__retimed_I5765_QOUT;
reg x_reg_L1_21__retimed_I5763_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5763_QOUT <= N10583;
	end
assign N10639 = x_reg_L1_21__retimed_I5763_QOUT;
reg x_reg_L1_21__retimed_I5762_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5762_QOUT <= N10581;
	end
assign N10637 = x_reg_L1_21__retimed_I5762_QOUT;
reg x_reg_L1_21__retimed_I5760_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5760_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3];
	end
assign N10632 = x_reg_L1_21__retimed_I5760_QOUT;
reg x_reg_L1_21__retimed_I5759_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5759_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7];
	end
assign N10630 = x_reg_L1_21__retimed_I5759_QOUT;
reg x_reg_L1_21__retimed_I5758_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5758_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5];
	end
assign N10627 = x_reg_L1_21__retimed_I5758_QOUT;
reg x_reg_L1_21__retimed_I5757_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5757_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4];
	end
assign N10625 = x_reg_L1_21__retimed_I5757_QOUT;
reg x_reg_L1_21__retimed_I5756_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5756_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2];
	end
assign N10623 = x_reg_L1_21__retimed_I5756_QOUT;
reg x_reg_L1_21__retimed_I5755_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5755_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0];
	end
assign N10621 = x_reg_L1_21__retimed_I5755_QOUT;
reg x_reg_L1_21__retimed_I5753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5753_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8];
	end
assign N10616 = x_reg_L1_21__retimed_I5753_QOUT;
reg x_reg_L0_21__retimed_I5739_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5739_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27;
	end
assign N10583 = x_reg_L0_21__retimed_I5739_QOUT;
reg x_reg_L0_21__retimed_I5738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5738_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28;
	end
assign N10581 = x_reg_L0_21__retimed_I5738_QOUT;
reg x_reg_L1_21__retimed_I5712_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5712_QOUT <= N9592;
	end
assign N10490 = x_reg_L1_21__retimed_I5712_QOUT;
reg x_reg_L1_21__retimed_I5710_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5710_QOUT <= N9566;
	end
assign N10464 = x_reg_L1_21__retimed_I5710_QOUT;
reg x_reg_L1_21__retimed_I5708_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5708_QOUT <= N9540;
	end
assign N10438 = x_reg_L1_21__retimed_I5708_QOUT;
reg x_reg_L1_21__retimed_I5706_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5706_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44;
	end
assign N10412 = x_reg_L1_21__retimed_I5706_QOUT;
reg x_reg_L1_21__retimed_I5658_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5658_QOUT <= N9279;
	end
assign N10262 = x_reg_L1_21__retimed_I5658_QOUT;
reg x_reg_L1_20__retimed_I5656_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5656_QOUT <= N9274;
	end
assign N10257 = x_reg_L1_20__retimed_I5656_QOUT;
reg x_reg_L1_19__retimed_I5654_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5654_QOUT <= N9269;
	end
assign N10252 = x_reg_L1_19__retimed_I5654_QOUT;
reg x_reg_L1_18__retimed_I5652_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5652_QOUT <= N9264;
	end
assign N10247 = x_reg_L1_18__retimed_I5652_QOUT;
reg x_reg_L1_17__retimed_I5650_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5650_QOUT <= N9259;
	end
assign N10242 = x_reg_L1_17__retimed_I5650_QOUT;
reg x_reg_L1_16__retimed_I5648_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5648_QOUT <= N9254;
	end
assign N10237 = x_reg_L1_16__retimed_I5648_QOUT;
reg x_reg_L1_15__retimed_I5646_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5646_QOUT <= N9249;
	end
assign N10232 = x_reg_L1_15__retimed_I5646_QOUT;
reg x_reg_L1_14__retimed_I5644_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5644_QOUT <= N9244;
	end
assign N10227 = x_reg_L1_14__retimed_I5644_QOUT;
reg x_reg_L1_13__retimed_I5642_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5642_QOUT <= N9239;
	end
assign N10222 = x_reg_L1_13__retimed_I5642_QOUT;
reg x_reg_L1_12__retimed_I5640_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5640_QOUT <= N9234;
	end
assign N10217 = x_reg_L1_12__retimed_I5640_QOUT;
reg x_reg_L1_11__retimed_I5638_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5638_QOUT <= N9229;
	end
assign N10212 = x_reg_L1_11__retimed_I5638_QOUT;
reg x_reg_L1_10__retimed_I5636_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5636_QOUT <= N9224;
	end
assign N10207 = x_reg_L1_10__retimed_I5636_QOUT;
reg x_reg_L1_9__retimed_I5634_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5634_QOUT <= N9219;
	end
assign N10202 = x_reg_L1_9__retimed_I5634_QOUT;
reg x_reg_L1_8__retimed_I5632_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5632_QOUT <= N9214;
	end
assign N10197 = x_reg_L1_8__retimed_I5632_QOUT;
reg x_reg_L1_7__retimed_I5630_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5630_QOUT <= N9209;
	end
assign N10192 = x_reg_L1_7__retimed_I5630_QOUT;
reg x_reg_L1_6__retimed_I5628_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5628_QOUT <= N9204;
	end
assign N10187 = x_reg_L1_6__retimed_I5628_QOUT;
reg x_reg_L1_5__retimed_I5626_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5626_QOUT <= N9199;
	end
assign N10182 = x_reg_L1_5__retimed_I5626_QOUT;
reg x_reg_L1_4__retimed_I5624_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5624_QOUT <= N9194;
	end
assign N10177 = x_reg_L1_4__retimed_I5624_QOUT;
reg x_reg_L1_3__retimed_I5622_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5622_QOUT <= N9189;
	end
assign N10172 = x_reg_L1_3__retimed_I5622_QOUT;
reg x_reg_L1_2__retimed_I5620_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5620_QOUT <= N9184;
	end
assign N10167 = x_reg_L1_2__retimed_I5620_QOUT;
reg x_reg_L1_1__retimed_I5618_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5618_QOUT <= N9179;
	end
assign N10162 = x_reg_L1_1__retimed_I5618_QOUT;
reg x_reg_L1_0__retimed_I5616_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5616_QOUT <= N9174;
	end
assign N10157 = x_reg_L1_0__retimed_I5616_QOUT;
reg x_reg_L1_21__retimed_I5614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5614_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45];
	end
assign N10152 = x_reg_L1_21__retimed_I5614_QOUT;
reg x_reg_L1_21__retimed_I5611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5611_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21];
	end
assign N10146 = x_reg_L1_21__retimed_I5611_QOUT;
reg x_reg_L1_20__retimed_I5610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5610_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44];
	end
assign N10143 = x_reg_L1_20__retimed_I5610_QOUT;
reg x_reg_L1_20__retimed_I5607_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5607_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20];
	end
assign N10137 = x_reg_L1_20__retimed_I5607_QOUT;
reg x_reg_L1_19__retimed_I5606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5606_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43];
	end
assign N10134 = x_reg_L1_19__retimed_I5606_QOUT;
reg x_reg_L1_19__retimed_I5603_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5603_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19];
	end
assign N10128 = x_reg_L1_19__retimed_I5603_QOUT;
reg x_reg_L1_18__retimed_I5602_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5602_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42];
	end
assign N10125 = x_reg_L1_18__retimed_I5602_QOUT;
reg x_reg_L1_18__retimed_I5599_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5599_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18];
	end
assign N10119 = x_reg_L1_18__retimed_I5599_QOUT;
reg x_reg_L1_17__retimed_I5598_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5598_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41];
	end
assign N10116 = x_reg_L1_17__retimed_I5598_QOUT;
reg x_reg_L1_17__retimed_I5595_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5595_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17];
	end
assign N10110 = x_reg_L1_17__retimed_I5595_QOUT;
reg x_reg_L1_16__retimed_I5594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5594_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40];
	end
assign N10107 = x_reg_L1_16__retimed_I5594_QOUT;
reg x_reg_L1_16__retimed_I5591_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5591_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16];
	end
assign N10101 = x_reg_L1_16__retimed_I5591_QOUT;
reg x_reg_L1_15__retimed_I5590_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5590_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39];
	end
assign N10098 = x_reg_L1_15__retimed_I5590_QOUT;
reg x_reg_L1_15__retimed_I5587_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5587_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15];
	end
assign N10092 = x_reg_L1_15__retimed_I5587_QOUT;
reg x_reg_L1_14__retimed_I5586_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5586_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38];
	end
assign N10089 = x_reg_L1_14__retimed_I5586_QOUT;
reg x_reg_L1_14__retimed_I5583_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5583_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14];
	end
assign N10083 = x_reg_L1_14__retimed_I5583_QOUT;
reg x_reg_L1_13__retimed_I5582_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5582_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37];
	end
assign N10080 = x_reg_L1_13__retimed_I5582_QOUT;
reg x_reg_L1_13__retimed_I5579_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5579_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13];
	end
assign N10074 = x_reg_L1_13__retimed_I5579_QOUT;
reg x_reg_L1_12__retimed_I5578_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5578_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36];
	end
assign N10071 = x_reg_L1_12__retimed_I5578_QOUT;
reg x_reg_L1_12__retimed_I5575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5575_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12];
	end
assign N10065 = x_reg_L1_12__retimed_I5575_QOUT;
reg x_reg_L1_11__retimed_I5574_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5574_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35];
	end
assign N10062 = x_reg_L1_11__retimed_I5574_QOUT;
reg x_reg_L1_11__retimed_I5571_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5571_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11];
	end
assign N10056 = x_reg_L1_11__retimed_I5571_QOUT;
reg x_reg_L1_10__retimed_I5570_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5570_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34];
	end
assign N10053 = x_reg_L1_10__retimed_I5570_QOUT;
reg x_reg_L1_10__retimed_I5567_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5567_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10];
	end
assign N10047 = x_reg_L1_10__retimed_I5567_QOUT;
reg x_reg_L1_9__retimed_I5566_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5566_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33];
	end
assign N10044 = x_reg_L1_9__retimed_I5566_QOUT;
reg x_reg_L1_9__retimed_I5563_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5563_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9];
	end
assign N10038 = x_reg_L1_9__retimed_I5563_QOUT;
reg x_reg_L1_8__retimed_I5562_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5562_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32];
	end
assign N10035 = x_reg_L1_8__retimed_I5562_QOUT;
reg x_reg_L1_8__retimed_I5559_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5559_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8];
	end
assign N10029 = x_reg_L1_8__retimed_I5559_QOUT;
reg x_reg_L1_7__retimed_I5558_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5558_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31];
	end
assign N10026 = x_reg_L1_7__retimed_I5558_QOUT;
reg x_reg_L1_7__retimed_I5555_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5555_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7];
	end
assign N10020 = x_reg_L1_7__retimed_I5555_QOUT;
reg x_reg_L1_6__retimed_I5554_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5554_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30];
	end
assign N10017 = x_reg_L1_6__retimed_I5554_QOUT;
reg x_reg_L1_6__retimed_I5551_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5551_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6];
	end
assign N10011 = x_reg_L1_6__retimed_I5551_QOUT;
reg x_reg_L1_5__retimed_I5550_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5550_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29];
	end
assign N10008 = x_reg_L1_5__retimed_I5550_QOUT;
reg x_reg_L1_5__retimed_I5547_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5547_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5];
	end
assign N10002 = x_reg_L1_5__retimed_I5547_QOUT;
reg x_reg_L1_4__retimed_I5546_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5546_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28];
	end
assign N9999 = x_reg_L1_4__retimed_I5546_QOUT;
reg x_reg_L1_4__retimed_I5543_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5543_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4];
	end
assign N9993 = x_reg_L1_4__retimed_I5543_QOUT;
reg x_reg_L1_3__retimed_I5542_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5542_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27];
	end
assign N9990 = x_reg_L1_3__retimed_I5542_QOUT;
reg x_reg_L1_3__retimed_I5539_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5539_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3];
	end
assign N9984 = x_reg_L1_3__retimed_I5539_QOUT;
reg x_reg_L1_2__retimed_I5538_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5538_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26];
	end
assign N9981 = x_reg_L1_2__retimed_I5538_QOUT;
reg x_reg_L1_2__retimed_I5535_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5535_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2];
	end
assign N9975 = x_reg_L1_2__retimed_I5535_QOUT;
reg x_reg_L1_1__retimed_I5534_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5534_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25];
	end
assign N9972 = x_reg_L1_1__retimed_I5534_QOUT;
reg x_reg_L1_1__retimed_I5531_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5531_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1];
	end
assign N9966 = x_reg_L1_1__retimed_I5531_QOUT;
reg x_reg_L1_0__retimed_I5530_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5530_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24];
	end
assign N9963 = x_reg_L1_0__retimed_I5530_QOUT;
reg x_reg_L1_0__retimed_I5527_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5527_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0];
	end
assign N9957 = x_reg_L1_0__retimed_I5527_QOUT;
reg x_reg_L1_21__retimed_I5523_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_21__retimed_I5523_QOUT <= N8965;
	end
assign N9948 = x_reg_L1_21__retimed_I5523_QOUT;
reg x_reg_L1_20__retimed_I5519_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_20__retimed_I5519_QOUT <= N8956;
	end
assign N9939 = x_reg_L1_20__retimed_I5519_QOUT;
reg x_reg_L1_19__retimed_I5515_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_19__retimed_I5515_QOUT <= N8947;
	end
assign N9930 = x_reg_L1_19__retimed_I5515_QOUT;
reg x_reg_L1_18__retimed_I5511_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_18__retimed_I5511_QOUT <= N8938;
	end
assign N9921 = x_reg_L1_18__retimed_I5511_QOUT;
reg x_reg_L1_17__retimed_I5507_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_17__retimed_I5507_QOUT <= N8929;
	end
assign N9912 = x_reg_L1_17__retimed_I5507_QOUT;
reg x_reg_L1_16__retimed_I5503_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_16__retimed_I5503_QOUT <= N8920;
	end
assign N9903 = x_reg_L1_16__retimed_I5503_QOUT;
reg x_reg_L1_15__retimed_I5499_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_15__retimed_I5499_QOUT <= N8911;
	end
assign N9894 = x_reg_L1_15__retimed_I5499_QOUT;
reg x_reg_L1_14__retimed_I5495_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_14__retimed_I5495_QOUT <= N8902;
	end
assign N9885 = x_reg_L1_14__retimed_I5495_QOUT;
reg x_reg_L1_13__retimed_I5491_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_13__retimed_I5491_QOUT <= N8893;
	end
assign N9876 = x_reg_L1_13__retimed_I5491_QOUT;
reg x_reg_L1_12__retimed_I5487_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_12__retimed_I5487_QOUT <= N8884;
	end
assign N9867 = x_reg_L1_12__retimed_I5487_QOUT;
reg x_reg_L1_11__retimed_I5483_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_11__retimed_I5483_QOUT <= N8875;
	end
assign N9858 = x_reg_L1_11__retimed_I5483_QOUT;
reg x_reg_L1_10__retimed_I5479_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_10__retimed_I5479_QOUT <= N8866;
	end
assign N9849 = x_reg_L1_10__retimed_I5479_QOUT;
reg x_reg_L1_9__retimed_I5475_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_9__retimed_I5475_QOUT <= N8857;
	end
assign N9840 = x_reg_L1_9__retimed_I5475_QOUT;
reg x_reg_L1_8__retimed_I5471_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_8__retimed_I5471_QOUT <= N8848;
	end
assign N9831 = x_reg_L1_8__retimed_I5471_QOUT;
reg x_reg_L1_7__retimed_I5467_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_7__retimed_I5467_QOUT <= N8839;
	end
assign N9822 = x_reg_L1_7__retimed_I5467_QOUT;
reg x_reg_L1_6__retimed_I5463_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_6__retimed_I5463_QOUT <= N8830;
	end
assign N9813 = x_reg_L1_6__retimed_I5463_QOUT;
reg x_reg_L1_5__retimed_I5459_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_5__retimed_I5459_QOUT <= N8821;
	end
assign N9804 = x_reg_L1_5__retimed_I5459_QOUT;
reg x_reg_L1_4__retimed_I5455_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_4__retimed_I5455_QOUT <= N8812;
	end
assign N9795 = x_reg_L1_4__retimed_I5455_QOUT;
reg x_reg_L1_3__retimed_I5451_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_3__retimed_I5451_QOUT <= N8803;
	end
assign N9786 = x_reg_L1_3__retimed_I5451_QOUT;
reg x_reg_L1_2__retimed_I5447_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_2__retimed_I5447_QOUT <= N8794;
	end
assign N9777 = x_reg_L1_2__retimed_I5447_QOUT;
reg x_reg_L1_1__retimed_I5443_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_1__retimed_I5443_QOUT <= N8785;
	end
assign N9768 = x_reg_L1_1__retimed_I5443_QOUT;
reg x_reg_L1_0__retimed_I5442_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5442_QOUT <= N8782;
	end
assign N9765 = x_reg_L1_0__retimed_I5442_QOUT;
assign N12999 = !N9765;
assign N13000 = !N12999;
reg x_reg_L1_0__retimed_I5439_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_0__retimed_I5439_QOUT <= N8776;
	end
assign N9759 = x_reg_L1_0__retimed_I5439_QOUT;
reg x_reg_L0_21__retimed_I5389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5389_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26;
	end
assign N9592 = x_reg_L0_21__retimed_I5389_QOUT;
reg x_reg_L0_21__retimed_I5387_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5387_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014;
	end
assign N9566 = x_reg_L0_21__retimed_I5387_QOUT;
reg x_reg_L0_21__retimed_I5385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5385_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095;
	end
assign N9540 = x_reg_L0_21__retimed_I5385_QOUT;
reg x_reg_L1_22__retimed_I5383_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5383_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923;
	end
assign N9514 = x_reg_L1_22__retimed_I5383_QOUT;
reg x_reg_L1_22__retimed_I5382_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_22__retimed_I5382_QOUT <= N8769;
	end
assign N9512 = x_reg_L1_22__retimed_I5382_QOUT;
reg x_reg_L1_23__retimed_I5380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5380_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870;
	end
assign N9507 = x_reg_L1_23__retimed_I5380_QOUT;
reg x_reg_L1_23__retimed_I5379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_23__retimed_I5379_QOUT <= N8762;
	end
assign N9505 = x_reg_L1_23__retimed_I5379_QOUT;
reg x_reg_L1_29__retimed_I5363_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_29__retimed_I5363_QOUT <= N8724;
	end
assign N9467 = x_reg_L1_29__retimed_I5363_QOUT;
reg x_reg_L0_21__retimed_I5286_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5286_QOUT <= a_man[21];
	end
assign N9279 = x_reg_L0_21__retimed_I5286_QOUT;
reg x_reg_L0_20__retimed_I5284_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5284_QOUT <= a_man[20];
	end
assign N9274 = x_reg_L0_20__retimed_I5284_QOUT;
reg x_reg_L0_19__retimed_I5282_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5282_QOUT <= a_man[19];
	end
assign N9269 = x_reg_L0_19__retimed_I5282_QOUT;
reg x_reg_L0_18__retimed_I5280_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5280_QOUT <= a_man[18];
	end
assign N9264 = x_reg_L0_18__retimed_I5280_QOUT;
reg x_reg_L0_17__retimed_I5278_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5278_QOUT <= a_man[17];
	end
assign N9259 = x_reg_L0_17__retimed_I5278_QOUT;
reg x_reg_L0_16__retimed_I5276_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5276_QOUT <= a_man[16];
	end
assign N9254 = x_reg_L0_16__retimed_I5276_QOUT;
reg x_reg_L0_15__retimed_I5274_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5274_QOUT <= a_man[15];
	end
assign N9249 = x_reg_L0_15__retimed_I5274_QOUT;
reg x_reg_L0_14__retimed_I5272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5272_QOUT <= a_man[14];
	end
assign N9244 = x_reg_L0_14__retimed_I5272_QOUT;
reg x_reg_L0_13__retimed_I5270_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5270_QOUT <= a_man[13];
	end
assign N9239 = x_reg_L0_13__retimed_I5270_QOUT;
reg x_reg_L0_12__retimed_I5268_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5268_QOUT <= a_man[12];
	end
assign N9234 = x_reg_L0_12__retimed_I5268_QOUT;
reg x_reg_L0_11__retimed_I5266_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5266_QOUT <= a_man[11];
	end
assign N9229 = x_reg_L0_11__retimed_I5266_QOUT;
reg x_reg_L0_10__retimed_I5264_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5264_QOUT <= a_man[10];
	end
assign N9224 = x_reg_L0_10__retimed_I5264_QOUT;
reg x_reg_L0_9__retimed_I5262_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5262_QOUT <= a_man[9];
	end
assign N9219 = x_reg_L0_9__retimed_I5262_QOUT;
reg x_reg_L0_8__retimed_I5260_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5260_QOUT <= a_man[8];
	end
assign N9214 = x_reg_L0_8__retimed_I5260_QOUT;
reg x_reg_L0_7__retimed_I5258_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5258_QOUT <= a_man[7];
	end
assign N9209 = x_reg_L0_7__retimed_I5258_QOUT;
reg x_reg_L0_6__retimed_I5256_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5256_QOUT <= a_man[6];
	end
assign N9204 = x_reg_L0_6__retimed_I5256_QOUT;
reg x_reg_L0_5__retimed_I5254_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5254_QOUT <= a_man[5];
	end
assign N9199 = x_reg_L0_5__retimed_I5254_QOUT;
reg x_reg_L0_4__retimed_I5252_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5252_QOUT <= a_man[4];
	end
assign N9194 = x_reg_L0_4__retimed_I5252_QOUT;
reg x_reg_L0_3__retimed_I5250_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5250_QOUT <= a_man[3];
	end
assign N9189 = x_reg_L0_3__retimed_I5250_QOUT;
reg x_reg_L0_2__retimed_I5248_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5248_QOUT <= a_man[2];
	end
assign N9184 = x_reg_L0_2__retimed_I5248_QOUT;
reg x_reg_L0_1__retimed_I5246_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5246_QOUT <= a_man[1];
	end
assign N9179 = x_reg_L0_1__retimed_I5246_QOUT;
reg x_reg_L0_0__retimed_I5244_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5244_QOUT <= a_man[0];
	end
assign N9174 = x_reg_L0_0__retimed_I5244_QOUT;
reg x_reg_L0_21__retimed_I5151_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_21__retimed_I5151_QOUT <= b_man[21];
	end
assign N8965 = x_reg_L0_21__retimed_I5151_QOUT;
reg x_reg_L0_20__retimed_I5147_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_20__retimed_I5147_QOUT <= b_man[20];
	end
assign N8956 = x_reg_L0_20__retimed_I5147_QOUT;
reg x_reg_L0_19__retimed_I5143_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_19__retimed_I5143_QOUT <= b_man[19];
	end
assign N8947 = x_reg_L0_19__retimed_I5143_QOUT;
reg x_reg_L0_18__retimed_I5139_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_18__retimed_I5139_QOUT <= b_man[18];
	end
assign N8938 = x_reg_L0_18__retimed_I5139_QOUT;
reg x_reg_L0_17__retimed_I5135_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_17__retimed_I5135_QOUT <= b_man[17];
	end
assign N8929 = x_reg_L0_17__retimed_I5135_QOUT;
reg x_reg_L0_16__retimed_I5131_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_16__retimed_I5131_QOUT <= b_man[16];
	end
assign N8920 = x_reg_L0_16__retimed_I5131_QOUT;
reg x_reg_L0_15__retimed_I5127_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_15__retimed_I5127_QOUT <= b_man[15];
	end
assign N8911 = x_reg_L0_15__retimed_I5127_QOUT;
reg x_reg_L0_14__retimed_I5123_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_14__retimed_I5123_QOUT <= b_man[14];
	end
assign N8902 = x_reg_L0_14__retimed_I5123_QOUT;
reg x_reg_L0_13__retimed_I5119_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_13__retimed_I5119_QOUT <= b_man[13];
	end
assign N8893 = x_reg_L0_13__retimed_I5119_QOUT;
reg x_reg_L0_12__retimed_I5115_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_12__retimed_I5115_QOUT <= b_man[12];
	end
assign N8884 = x_reg_L0_12__retimed_I5115_QOUT;
reg x_reg_L0_11__retimed_I5111_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_11__retimed_I5111_QOUT <= b_man[11];
	end
assign N8875 = x_reg_L0_11__retimed_I5111_QOUT;
reg x_reg_L0_10__retimed_I5107_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_10__retimed_I5107_QOUT <= b_man[10];
	end
assign N8866 = x_reg_L0_10__retimed_I5107_QOUT;
reg x_reg_L0_9__retimed_I5103_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_9__retimed_I5103_QOUT <= b_man[9];
	end
assign N8857 = x_reg_L0_9__retimed_I5103_QOUT;
reg x_reg_L0_8__retimed_I5099_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_8__retimed_I5099_QOUT <= b_man[8];
	end
assign N8848 = x_reg_L0_8__retimed_I5099_QOUT;
reg x_reg_L0_7__retimed_I5095_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_7__retimed_I5095_QOUT <= b_man[7];
	end
assign N8839 = x_reg_L0_7__retimed_I5095_QOUT;
reg x_reg_L0_6__retimed_I5091_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_6__retimed_I5091_QOUT <= b_man[6];
	end
assign N8830 = x_reg_L0_6__retimed_I5091_QOUT;
reg x_reg_L0_5__retimed_I5087_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_5__retimed_I5087_QOUT <= b_man[5];
	end
assign N8821 = x_reg_L0_5__retimed_I5087_QOUT;
reg x_reg_L0_4__retimed_I5083_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_4__retimed_I5083_QOUT <= b_man[4];
	end
assign N8812 = x_reg_L0_4__retimed_I5083_QOUT;
reg x_reg_L0_3__retimed_I5079_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_3__retimed_I5079_QOUT <= b_man[3];
	end
assign N8803 = x_reg_L0_3__retimed_I5079_QOUT;
reg x_reg_L0_2__retimed_I5075_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_2__retimed_I5075_QOUT <= b_man[2];
	end
assign N8794 = x_reg_L0_2__retimed_I5075_QOUT;
reg x_reg_L0_1__retimed_I5071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_1__retimed_I5071_QOUT <= b_man[1];
	end
assign N8785 = x_reg_L0_1__retimed_I5071_QOUT;
reg x_reg_L0_0__retimed_I5070_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5070_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47;
	end
assign N8782 = x_reg_L0_0__retimed_I5070_QOUT;
reg x_reg_L0_0__retimed_I5067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_0__retimed_I5067_QOUT <= b_man[0];
	end
assign N8776 = x_reg_L0_0__retimed_I5067_QOUT;
reg x_reg_L0_22__retimed_I5064_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_22__retimed_I5064_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925;
	end
assign N8769 = x_reg_L0_22__retimed_I5064_QOUT;
reg x_reg_L0_23__retimed_I5061_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_23__retimed_I5061_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893;
	end
assign N8762 = x_reg_L0_23__retimed_I5061_QOUT;
reg x_reg_L0_29__retimed_I5045_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_29__retimed_I5045_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874;
	end
assign N8724 = x_reg_L0_29__retimed_I5045_QOUT;
assign bdw_enable = !astall;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011 = !(a_exp[0] & a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013 = ((a_exp[5] & a_exp[4]) & a_exp[3]) & a_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396 = !((a_exp[7] & a_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047 = ((a_man[22] | a_man[20]) | a_man[21]) | a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051 = !(((a_man[0] | a_man[1]) | a_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034 = !(a_man[10] | a_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053 = !(a_man[6] | a_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042 = !(a_man[8] | a_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062 = !(a_man[4] | a_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056 = ((a_man[18] | a_man[16]) | a_man[17]) | a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066 = ((a_man[14] | a_man[12]) | a_man[13]) | a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900 = !(b_exp[0] & b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902 = ((b_exp[5] & b_exp[4]) & b_exp[3]) & b_exp[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388 = !((b_exp[7] & b_exp[6]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936 = ((b_man[22] | b_man[20]) | b_man[21]) | b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940 = !(((b_man[0] | b_man[1]) | b_man[2]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923 = !(b_man[10] | b_man[9]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942 = !(b_man[6] | b_man[5]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931 = !(b_man[8] | b_man[7]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951 = !(b_man[4] | b_man[3]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945 = ((b_man[18] | b_man[16]) | b_man[17]) | b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955 = ((b_man[14] | b_man[12]) | b_man[13]) | b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985 = !(a_exp[0] | a_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992 = !(a_exp[5] | a_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989 = !(a_exp[7] | a_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980 = !(a_exp[3] | a_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096 = !(b_exp[0] | b_exp[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103 = !(b_exp[5] | b_exp[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100 = !(b_exp[7] | b_exp[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091 = !(b_exp[3] | b_exp[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0] = (!b_exp[0]) ^ a_exp[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134 = !a_man[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320 = (!b_man[22]) ^ b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452 = !a_man[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799 = !a_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963 = b_man[22] | b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385 = (!b_man[20]) ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118 = b_man[21] ^ b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395 = !b_man[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329 = !a_man[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660 = !a_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450 = (!b_man[18]) ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325 = b_man[19] ^ b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993 = !b_man[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653 = !a_man[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987 = !a_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090 = b_man[17] ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519 = (!b_man[16]) ^ b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583 = !b_man[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513 = !a_man[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308 = !a_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586 = (!b_man[14]) ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295 = b_man[15] ^ b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352 = !b_man[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853 = !a_man[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186 = !a_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646 = (!b_man[12]) ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060 = b_man[13] ^ b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947 = !b_man[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171 = !a_man[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511 = !a_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712 = (!b_man[10]) ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267 = b_man[11] ^ b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258 = !b_man[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047 = !a_man[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391 = !a_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779 = (!b_man[8]) ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033 = b_man[9] ^ b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564 = !b_man[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368 = !a_man[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713 = !a_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844 = (!b_man[6]) ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242 = b_man[7] ^ b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332 = !b_man[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243 = !a_man[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578 = !a_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906 = b_man[4] ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004 = (!b_man[5]) ^ b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645 = !b_man[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573 = !a_man[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911 = !a_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968 = (!b_man[2]) ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211 = b_man[3] ^ b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959 = !b_man[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228 = !a_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445 = !a_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272 = !b_man[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357 = !b_man[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935 = !(b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807 = !(b_man[21] & b_man[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529 = !(b_man[19] & b_man[20]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871 = b_man[21] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595 = !(b_man[17] & b_man[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933 = b_man[19] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658 = !(b_man[15] & b_man[16]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994 = b_man[17] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721 = !(b_man[13] & b_man[14]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058 = b_man[15] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795 = !(b_man[11] & b_man[12]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126 = b_man[13] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855 = !(b_man[9] & b_man[10]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185 = b_man[11] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916 = !(b_man[7] & b_man[8]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251 = b_man[9] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978 = !(b_man[5] & b_man[6]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317 = b_man[7] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045 = !(b_man[3] & b_man[4]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385 = b_man[5] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913};
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111 = !(b_man[1] & b_man[2]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446 = b_man[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290} = {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357)) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435 = b_man[1] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558) & (!(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922) & (!(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728)));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151 = (!N11830) | (N11566 & N11564);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393 = (!N11822) | (N11560 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197 = (!N11814) | (N11554 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239 = (!N11806) | (N11548 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412 = (!N11798) | (N11542 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701 = (!N11790) | (N11536 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670 = (!N11782) | (N11530 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310 = (!N11774) | (N11524 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081 = (!N11766) | (N11518 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516 = (!N11758) | (N11512 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104 = (!N11750) | (N11506 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349 = (!N11742) | (N11500 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723 = (!N11734) | (N11177 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776 = (!N11726) | (N11171 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493 = (!N11718) | (N11165 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356 = (!N11710) | (N11159 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331 = (!N11702) | (N11153 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526 = (!N11694) | (N11147 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315 = (!N11686) | (N11141 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326 = (!N11678) | (N11135 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326 ^ N11675;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315) ^ N11135;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356) ^ N11153;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331) ^ N11147;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493) ^ N11159;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526) ^ N11141;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393) ^ N11554;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197) ^ N11548;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151) ^ N11560;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27] = (!N11564) ^ N11566;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26] = (!N11570) ^ N11572;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11241);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11241) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11239);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11239) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10847);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0] = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516) ^ N11506;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104) ^ N11500;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081) ^ N11512;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310) ^ N11518;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670) ^ N11524;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701) ^ N11530;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412) ^ N11536;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239) ^ N11542;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776) ^ N11165;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723) ^ N11171;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349) ^ N11177;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24] = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10847) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N10845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8 = !(((!rm[2]) | rm[1]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 = !(((!rm[1]) | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23 = a_sign ^ b_sign;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 = !(((!rm[0]) | rm[2]) | rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11366) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11364);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11387) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11385);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11408) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11406);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11345) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11343);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11352) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11350);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11373) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11359);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11357) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11378) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11401);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11359) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11357);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11364) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11378);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11401) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11406) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11366);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11392) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11352);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N10845) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11449);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11447) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11454);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224 = ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11470) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11468);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0] = b_man[1] ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11475;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376 & N11350) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376) & N11475);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373 & N11449) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373) & N11447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N11454) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N11470);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N11468) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N11345);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N11343) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N11387);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224 & N11385) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224) & N11408);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4 = !((rm[1] | rm[2]) | rm[0]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24])) | (!N10872));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447 = ((N10827 | N10829) | N10831) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450 = ((!N10831) & (!N10829)) | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10696) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10694);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631 = b_exp[0] | a_exp[0];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]} = {1'B0, a_exp[1]} + {1'B0, b_exp[1]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0] | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]));
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]} = {1'B0, a_exp[2]} + {1'B0, b_exp[2]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10705) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10703);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]} = {1'B0, a_exp[3]} + {1'B0, b_exp[3]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682;
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]} = {1'B0, a_exp[4]} + {1'B0, b_exp[4]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10714) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10712);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]} = {1'B0, a_exp[5]} + {1'B0, b_exp[5]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10723) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10721);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812 = !(((N10621 | N10623) | N10625) | N10627);
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]} = {1'B0, a_exp[6]} + {1'B0, b_exp[6]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627 = !a_exp[7];
assign {float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]} = {1'B0, b_exp[7]} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627} + {1'B0, float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632};
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10741) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10739);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10759) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10757);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] = (!a_exp[7]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10776) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10774);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10768) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10766);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813 = !(N10616 | N11432);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10750) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10748);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9] = !(a_exp[7] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38 & N10732) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38) & N10730);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801 = !(N11425 | N10643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808 = !((N10630 | N10632) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830 = !(((N10637 | N10639) | N10490) | N10643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823 = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768 = !(N11432 & N11425);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763 = !(N10630 & N10632);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775 = !(N10625 & N10623);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772 = !(N10621 & N10627);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461 = !(((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417 = !(N10616 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417 | N10643);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 = !(N10438 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10262);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028 = N10412 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887;
assign N13001 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028;
assign N13002 = !N13001;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 = !(N10412 | (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951 = !((N13002 & N10146) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10152));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380 = !(N10464 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign N13003 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380;
assign N13004 = !N13003;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 = !(N10490 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852 = !(rm[0] & rm[1]);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7 = !(rm[2] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914 = ((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8] | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043 = !((N13004 & N9948) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[21] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10257);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061 = !((N13002 & N10137) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10143));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069 = !((N13004 & N9939) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[20] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10252);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977 = !((N13002 & N10128) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10134));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091 = !((N13004 & N9930) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[19] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10247);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084 = !((N13002 & N10119) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10125));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117 = !((N13004 & N9921) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[18] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10242);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002 = !((N13002 & N10110) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10116));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948 = !((N13004 & N9912) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[17] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10237);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109 = !((N13002 & N10101) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10107));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973 = !((N13004 & N9903) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[16] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10232);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027 = !((N13002 & N10092) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10098));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999 = !((N13004 & N9894) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[15] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10227);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941 = !((N13002 & N10083) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10089));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024 = !((N13004 & N9885) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[14] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10222);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051 = !((N13002 & N10074) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10080));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047 = !((N13004 & N9876) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[13] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10217);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967 = !((N13002 & N10065) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10071));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073 = !((N13004 & N9867) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[12] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10212);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077 = !((N13002 & N10056) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10062));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096 = !((N13004 & N9858) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[11] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10207);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363 = !(((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992 = !((N13002 & N10047) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10053));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930 = !((N13004 & N9849) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[10] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10202);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100 = !((N13002 & N10038) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10044));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953 = !((N13004 & N9840) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[9] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10197);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018 = !((N13002 & N10029) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10035));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978 = !((N13004 & N9831) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[8] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10192);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933 = !((N13002 & N10020) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10026));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004 = !((N13004 & N9822) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[7] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10187);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]) & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040 = !((N13002 & N10011) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10017));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030 = !((N13004 & N9813) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[6] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10182);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957 = !((N13002 & N10002) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N10008));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053 = !((N13004 & N9804) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[5] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10177);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27] & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066 = !((N13002 & N9993) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N9999));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079 = !((N13004 & N9795) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[4] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10172);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3] = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387 ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982 = !((N13002 & N9984) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N9990));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102 = !((N13004 & N9786) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[3] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10167);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25] & (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088 = !((N13002 & N9975) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N9981));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934 = !((N13004 & N9777) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[2] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10162);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008 = !((N13002 & N9966) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N9972));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959 = !((N13004 & N9768) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[1] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382 & N10157);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114 = !((N13002 & N9957) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987 & N9963));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984 = !((N13004 & N9759) | (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378 & N13000));
assign x[0] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336 = !((((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22] = (!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336) ^ float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22]) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47);
assign x[22] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49 & N9512) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49) & N9514));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874 = float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887;
assign x[30] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N10630);
assign x[29] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N11425);
assign x[28] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N10627);
assign x[27] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N10625);
assign x[26] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N10632);
assign x[25] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N10623);
assign x[24] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9467) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N11432);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870 = !float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893 = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42) | float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470);
assign x[23] = !((float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884 & N9505) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884) & N9507));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135 = !(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22 & (!b_sign));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140 = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15 & a_sign) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135);
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31] = (float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26 & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140) | ((!float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26) & float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23);
reg x_reg_L0_31__I1625_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L0_31__I1625_QOUT <= float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31];
	end
assign N4032 = x_reg_L0_31__I1625_QOUT;
reg x_reg_L1_31__I1657_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_L1_31__I1657_QOUT <= N4032;
	end
assign x[31] = x_reg_L1_31__I1657_QOUT;
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vbD5SgzWrxA= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



