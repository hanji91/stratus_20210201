/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:28 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_mul_ieee_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable;
wire [31:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23;
wire [47:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44;
wire [24:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47;
wire [9:0] float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48;
wire  float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411,
	float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417;
wire N4032,N8724,N8762,N8769,N8776,N8782,N8785 
	,N8794,N8803,N8812,N8821,N8830,N8839,N8848,N8857 
	,N8866,N8875,N8884,N8893,N8902,N8911,N8920,N8929 
	,N8938,N8947,N8956,N8965,N9174,N9179,N9184,N9189 
	,N9194,N9199,N9204,N9209,N9214,N9219,N9224,N9229 
	,N9234,N9239,N9244,N9249,N9254,N9259,N9264,N9269 
	,N9274,N9279,N9467,N9505,N9507,N9512,N9514,N9540 
	,N9566,N9592,N9759,N9765,N9768,N9777,N9786,N9795 
	,N9804,N9813,N9822,N9831,N9840,N9849,N9858,N9867 
	,N9876,N9885,N9894,N9903,N9912,N9921,N9930,N9939 
	,N9948,N9957,N9963,N9966,N9972,N9975,N9981,N9984 
	,N9990,N9993,N9999,N10002,N10008,N10011,N10017,N10020 
	,N10026,N10029,N10035,N10038,N10044,N10047,N10053,N10056 
	,N10062,N10065,N10071,N10074,N10080,N10083,N10089,N10092 
	,N10098,N10101,N10107,N10110,N10116,N10119,N10125,N10128 
	,N10134,N10137,N10143,N10146,N10152,N10157,N10162,N10167 
	,N10172,N10177,N10182,N10187,N10192,N10197,N10202,N10207 
	,N10212,N10217,N10222,N10227,N10232,N10237,N10242,N10247 
	,N10252,N10257,N10262,N10412,N10438,N10464,N10490,N10581 
	,N10583,N10616,N10621,N10623,N10625,N10627,N10630,N10632 
	,N10637,N10639,N10643,N10694,N10696,N10703,N10705,N10712 
	,N10714,N10721,N10723,N10730,N10732,N10739,N10741,N10748 
	,N10750,N10757,N10759,N10766,N10768,N10774,N10776,N10827 
	,N10829,N10831,N10845,N10847,N10872,N11135,N11141,N11147 
	,N11153,N11159,N11165,N11171,N11177,N11239,N11241,N11343 
	,N11345,N11350,N11352,N11357,N11359,N11364,N11366,N11373 
	,N11378,N11385,N11387,N11392,N11401,N11406,N11408,N11425 
	,N11432,N11447,N11449,N11454,N11468,N11470,N11475,N11500 
	,N11506,N11512,N11518,N11524,N11530,N11536,N11542,N11548 
	,N11554,N11560,N11564,N11566,N11570,N11572,N11675,N11678 
	,N11686,N11694,N11702,N11710,N11718,N11726,N11734,N11742 
	,N11750,N11758,N11766,N11774,N11782,N11790,N11798,N11806 
	,N11814,N11822,N11830,N12999,N13000,N13001,N13002,N13003 
	,N13004;
EDFFHQX1 x_reg_L0_21__retimed_I6170 (.Q(N11830), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6167 (.Q(N11822), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6164 (.Q(N11814), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6161 (.Q(N11806), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6158 (.Q(N11798), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6155 (.Q(N11790), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6152 (.Q(N11782), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6149 (.Q(N11774), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6146 (.Q(N11766), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6143 (.Q(N11758), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6140 (.Q(N11750), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6137 (.Q(N11742), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6134 (.Q(N11734), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6131 (.Q(N11726), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6128 (.Q(N11718), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6125 (.Q(N11710), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6122 (.Q(N11702), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6119 (.Q(N11694), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6116 (.Q(N11686), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6113 (.Q(N11678), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6112 (.Q(N11675), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6090 (.Q(N11572), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6089 (.Q(N11570), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6088 (.Q(N11566), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6087 (.Q(N11564), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6086 (.Q(N11560), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6084 (.Q(N11554), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6082 (.Q(N11548), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6080 (.Q(N11542), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6078 (.Q(N11536), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6076 (.Q(N11530), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6074 (.Q(N11524), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6072 (.Q(N11518), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6070 (.Q(N11512), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6068 (.Q(N11506), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6066 (.Q(N11500), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6056 (.Q(N11475), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6054 (.Q(N11470), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6053 (.Q(N11468), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6047 (.Q(N11454), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6045 (.Q(N11449), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6044 (.Q(N11447), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I6038 (.Q(N11432), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I6035 (.Q(N11425), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6028 (.Q(N11408), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6027 (.Q(N11406), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6025 (.Q(N11401), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6021 (.Q(N11392), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6019 (.Q(N11387), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6018 (.Q(N11385), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6015 (.Q(N11378), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6013 (.Q(N11373), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6010 (.Q(N11366), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6009 (.Q(N11364), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6007 (.Q(N11359), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6006 (.Q(N11357), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6004 (.Q(N11352), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6003 (.Q(N11350), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6001 (.Q(N11345), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I6000 (.Q(N11343), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5966 (.Q(N11241), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5965 (.Q(N11239), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5945 (.Q(N11177), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5943 (.Q(N11171), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5941 (.Q(N11165), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5939 (.Q(N11159), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5937 (.Q(N11153), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5935 (.Q(N11147), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5933 (.Q(N11141), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5931 (.Q(N11135), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5845 (.Q(N10872), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5838 (.Q(N10847), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5837 (.Q(N10845), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5831 (.Q(N10831), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5830 (.Q(N10829), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5829 (.Q(N10827), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5813 (.Q(N10776), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5812 (.Q(N10774), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5810 (.Q(N10768), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5809 (.Q(N10766), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5807 (.Q(N10759), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5806 (.Q(N10757), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5804 (.Q(N10750), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5803 (.Q(N10748), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5801 (.Q(N10741), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5800 (.Q(N10739), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5798 (.Q(N10732), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5797 (.Q(N10730), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5795 (.Q(N10723), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5794 (.Q(N10721), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5792 (.Q(N10714), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5791 (.Q(N10712), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5789 (.Q(N10705), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5788 (.Q(N10703), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5786 (.Q(N10696), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5785 (.Q(N10694), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5765 (.Q(N10643), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5763 (.Q(N10639), .D(N10583), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5762 (.Q(N10637), .D(N10581), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5760 (.Q(N10632), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5759 (.Q(N10630), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5758 (.Q(N10627), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5757 (.Q(N10625), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5756 (.Q(N10623), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5755 (.Q(N10621), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5753 (.Q(N10616), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5739 (.Q(N10583), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5738 (.Q(N10581), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5712 (.Q(N10490), .D(N9592), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5710 (.Q(N10464), .D(N9566), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5708 (.Q(N10438), .D(N9540), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5706 (.Q(N10412), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5658 (.Q(N10262), .D(N9279), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I5656 (.Q(N10257), .D(N9274), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I5654 (.Q(N10252), .D(N9269), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I5652 (.Q(N10247), .D(N9264), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I5650 (.Q(N10242), .D(N9259), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I5648 (.Q(N10237), .D(N9254), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I5646 (.Q(N10232), .D(N9249), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I5644 (.Q(N10227), .D(N9244), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I5642 (.Q(N10222), .D(N9239), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I5640 (.Q(N10217), .D(N9234), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I5638 (.Q(N10212), .D(N9229), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I5636 (.Q(N10207), .D(N9224), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I5634 (.Q(N10202), .D(N9219), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I5632 (.Q(N10197), .D(N9214), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I5630 (.Q(N10192), .D(N9209), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I5628 (.Q(N10187), .D(N9204), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I5626 (.Q(N10182), .D(N9199), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I5624 (.Q(N10177), .D(N9194), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I5622 (.Q(N10172), .D(N9189), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I5620 (.Q(N10167), .D(N9184), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I5618 (.Q(N10162), .D(N9179), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I5616 (.Q(N10157), .D(N9174), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5614 (.Q(N10152), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5611 (.Q(N10146), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I5610 (.Q(N10143), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I5607 (.Q(N10137), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I5606 (.Q(N10134), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I5603 (.Q(N10128), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I5602 (.Q(N10125), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I5599 (.Q(N10119), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I5598 (.Q(N10116), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I5595 (.Q(N10110), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I5594 (.Q(N10107), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I5591 (.Q(N10101), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I5590 (.Q(N10098), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I5587 (.Q(N10092), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I5586 (.Q(N10089), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I5583 (.Q(N10083), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I5582 (.Q(N10080), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I5579 (.Q(N10074), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I5578 (.Q(N10071), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I5575 (.Q(N10065), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I5574 (.Q(N10062), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I5571 (.Q(N10056), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I5570 (.Q(N10053), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I5567 (.Q(N10047), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I5566 (.Q(N10044), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I5563 (.Q(N10038), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I5562 (.Q(N10035), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I5559 (.Q(N10029), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I5558 (.Q(N10026), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I5555 (.Q(N10020), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I5554 (.Q(N10017), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I5551 (.Q(N10011), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I5550 (.Q(N10008), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I5547 (.Q(N10002), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I5546 (.Q(N9999), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I5543 (.Q(N9993), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I5542 (.Q(N9990), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I5539 (.Q(N9984), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I5538 (.Q(N9981), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I5535 (.Q(N9975), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I5534 (.Q(N9972), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I5531 (.Q(N9966), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I5530 (.Q(N9963), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I5527 (.Q(N9957), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_21__retimed_I5523 (.Q(N9948), .D(N8965), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_20__retimed_I5519 (.Q(N9939), .D(N8956), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_19__retimed_I5515 (.Q(N9930), .D(N8947), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_18__retimed_I5511 (.Q(N9921), .D(N8938), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_17__retimed_I5507 (.Q(N9912), .D(N8929), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_16__retimed_I5503 (.Q(N9903), .D(N8920), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_15__retimed_I5499 (.Q(N9894), .D(N8911), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_14__retimed_I5495 (.Q(N9885), .D(N8902), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_13__retimed_I5491 (.Q(N9876), .D(N8893), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_12__retimed_I5487 (.Q(N9867), .D(N8884), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_11__retimed_I5483 (.Q(N9858), .D(N8875), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_10__retimed_I5479 (.Q(N9849), .D(N8866), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_9__retimed_I5475 (.Q(N9840), .D(N8857), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_8__retimed_I5471 (.Q(N9831), .D(N8848), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_7__retimed_I5467 (.Q(N9822), .D(N8839), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_6__retimed_I5463 (.Q(N9813), .D(N8830), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_5__retimed_I5459 (.Q(N9804), .D(N8821), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_4__retimed_I5455 (.Q(N9795), .D(N8812), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_3__retimed_I5451 (.Q(N9786), .D(N8803), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_2__retimed_I5447 (.Q(N9777), .D(N8794), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_1__retimed_I5443 (.Q(N9768), .D(N8785), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_0__retimed_I5442 (.Q(N9765), .D(N8782), .E(bdw_enable), .CK(aclk));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6693 (.Y(N12999), .A(N9765));
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6694 (.Y(N13000), .A(N12999));
EDFFHQX1 x_reg_L1_0__retimed_I5439 (.Q(N9759), .D(N8776), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5389 (.Q(N9592), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5387 (.Q(N9566), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5385 (.Q(N9540), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I5383 (.Q(N9514), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_22__retimed_I5382 (.Q(N9512), .D(N8769), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I5380 (.Q(N9507), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_23__retimed_I5379 (.Q(N9505), .D(N8762), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_29__retimed_I5363 (.Q(N9467), .D(N8724), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5286 (.Q(N9279), .D(a_man[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_20__retimed_I5284 (.Q(N9274), .D(a_man[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_19__retimed_I5282 (.Q(N9269), .D(a_man[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_18__retimed_I5280 (.Q(N9264), .D(a_man[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_17__retimed_I5278 (.Q(N9259), .D(a_man[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_16__retimed_I5276 (.Q(N9254), .D(a_man[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_15__retimed_I5274 (.Q(N9249), .D(a_man[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_14__retimed_I5272 (.Q(N9244), .D(a_man[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_13__retimed_I5270 (.Q(N9239), .D(a_man[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_12__retimed_I5268 (.Q(N9234), .D(a_man[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_11__retimed_I5266 (.Q(N9229), .D(a_man[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_10__retimed_I5264 (.Q(N9224), .D(a_man[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_9__retimed_I5262 (.Q(N9219), .D(a_man[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_8__retimed_I5260 (.Q(N9214), .D(a_man[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_7__retimed_I5258 (.Q(N9209), .D(a_man[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_6__retimed_I5256 (.Q(N9204), .D(a_man[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_5__retimed_I5254 (.Q(N9199), .D(a_man[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_4__retimed_I5252 (.Q(N9194), .D(a_man[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_3__retimed_I5250 (.Q(N9189), .D(a_man[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_2__retimed_I5248 (.Q(N9184), .D(a_man[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_1__retimed_I5246 (.Q(N9179), .D(a_man[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I5244 (.Q(N9174), .D(a_man[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_21__retimed_I5151 (.Q(N8965), .D(b_man[21]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_20__retimed_I5147 (.Q(N8956), .D(b_man[20]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_19__retimed_I5143 (.Q(N8947), .D(b_man[19]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_18__retimed_I5139 (.Q(N8938), .D(b_man[18]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_17__retimed_I5135 (.Q(N8929), .D(b_man[17]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_16__retimed_I5131 (.Q(N8920), .D(b_man[16]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_15__retimed_I5127 (.Q(N8911), .D(b_man[15]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_14__retimed_I5123 (.Q(N8902), .D(b_man[14]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_13__retimed_I5119 (.Q(N8893), .D(b_man[13]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_12__retimed_I5115 (.Q(N8884), .D(b_man[12]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_11__retimed_I5111 (.Q(N8875), .D(b_man[11]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_10__retimed_I5107 (.Q(N8866), .D(b_man[10]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_9__retimed_I5103 (.Q(N8857), .D(b_man[9]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_8__retimed_I5099 (.Q(N8848), .D(b_man[8]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_7__retimed_I5095 (.Q(N8839), .D(b_man[7]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_6__retimed_I5091 (.Q(N8830), .D(b_man[6]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_5__retimed_I5087 (.Q(N8821), .D(b_man[5]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_4__retimed_I5083 (.Q(N8812), .D(b_man[4]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_3__retimed_I5079 (.Q(N8803), .D(b_man[3]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_2__retimed_I5075 (.Q(N8794), .D(b_man[2]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_1__retimed_I5071 (.Q(N8785), .D(b_man[1]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I5070 (.Q(N8782), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_0__retimed_I5067 (.Q(N8776), .D(b_man[0]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_22__retimed_I5064 (.Q(N8769), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_23__retimed_I5061 (.Q(N8762), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L0_29__retimed_I5045 (.Q(N8724), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874), .E(bdw_enable), .CK(aclk));
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011), .A(a_exp[0]), .B(a_exp[1]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I2 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I3 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396), .A(a_exp[7]), .B(a_exp[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2013));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I4 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2011), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8396));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I5 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2047));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I7 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034), .A(a_man[10]), .B(a_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I8 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053), .A(a_man[6]), .B(a_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I9 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042), .A(a_man[8]), .B(a_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I10 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062), .A(a_man[4]), .B(a_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I11 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2034), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2053), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2042), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2062));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I12 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I13 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I14 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2051), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2045), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2056), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2066));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I15 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I16 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900), .A(b_exp[0]), .B(b_exp[1]));
AND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I17 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I18 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388), .A(b_exp[7]), .B(b_exp[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1902));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I19 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1900), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8388));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I20 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I21 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1936));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I22 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923), .A(b_man[10]), .B(b_man[9]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I23 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942), .A(b_man[6]), .B(b_man[5]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I24 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931), .A(b_man[8]), .B(b_man[7]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I25 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951), .A(b_man[4]), .B(b_man[3]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I26 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1923), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1942), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1931), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1951));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I27 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I28 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I29 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1940), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1934), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1945), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1955));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I30 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I31 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I32 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I33 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I34 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I35 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1985), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1992), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1989), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N1980));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I36 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__17), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__19));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I37 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I38 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096), .A(b_exp[0]), .B(b_exp[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I39 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103), .A(b_exp[5]), .B(b_exp[4]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I40 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100), .A(b_exp[7]), .B(b_exp[6]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I41 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091), .A(b_exp[3]), .B(b_exp[2]));
NAND4XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I42 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2096), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2103), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2100), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2091));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I43 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__10), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__12));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I44 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I45 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N441), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N440));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I46 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6095), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I47 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0]), .A(b_exp[0]), .B(a_exp[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I48 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I49 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .A(a_man[22]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I50 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .A(b_man[22]), .B(b_man[21]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I51 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I52 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .A(a_man[20]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I53 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I54 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .A(a_man[21]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I55 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I56 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I57 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963), .A(b_man[22]), .B(b_man[21]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I58 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I59 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2454));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I60 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3136), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3011));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I61 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .A(b_man[20]), .B(b_man[19]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I62 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118), .A(b_man[21]), .B(b_man[19]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I63 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3118), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I64 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395), .A(b_man[21]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I65 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I66 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I67 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I68 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3664), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I69 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I70 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2377), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3333), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2430));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I71 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2676), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2955), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3068));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I72 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2503), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I73 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .A(a_man[18]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I74 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I75 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .A(a_man[19]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I76 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I77 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2990), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I78 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2657));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I79 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .A(b_man[18]), .B(b_man[17]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I80 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325), .A(b_man[19]), .B(b_man[17]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I81 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2325), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I82 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993), .A(b_man[19]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I83 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I84 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I85 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3587), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I86 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2615), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3256), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2797));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I87 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2732), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3130), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3269));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I88 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3379), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I89 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I90 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2919), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I91 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2313), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I92 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I93 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2583), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3518), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2488));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I94 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .A(a_man[16]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I95 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I96 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .A(a_man[17]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I97 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I98 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3190), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I99 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2857));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I101 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I102 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2568), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2442), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2167));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I103 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2506), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3325));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I104 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2704), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I105 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I107 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2516), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I110 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2642), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2175), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3055));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2238), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090), .A(b_man[17]), .B(b_man[15]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .A(b_man[16]), .B(b_man[15]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I115 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3090), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I116 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583), .A(b_man[17]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I117 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I118 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I119 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3115), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .A(a_man[14]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I122 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .A(a_man[15]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3395), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I126 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3050));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I127 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2509), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2783), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2881));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I128 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2283), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3451), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3634));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I129 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3652), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2979), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I131 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3321), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2273), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2945));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I132 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2709), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2224), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2983));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I133 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3571), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I135 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2300), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I136 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I137 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2169), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2436), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I140 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3507), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3390), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3646));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I141 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3489), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2344), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3299));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I142 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2366), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3442), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3105));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I143 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2900), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I144 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586), .A(b_man[14]), .B(b_man[13]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I145 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I146 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I147 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295), .A(b_man[15]), .B(b_man[13]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2295), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2586));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I149 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352), .A(b_man[15]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .A(a_man[12]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I152 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .A(a_man[13]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I154 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I155 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I156 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3245));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I157 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I158 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I160 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I162 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I164 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I165 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I166 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2163), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3576), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2294));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I169 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3177), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2502), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I170 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3314), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2635), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I171 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2580), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2847), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2974));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I172 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3189), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2656), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2212));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I173 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2542), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3481), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2599));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3046), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2367), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I175 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2714), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3581), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I177 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2710), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2372), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3623));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I178 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2940), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2801), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3503));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I179 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2480), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3546), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3197));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2219), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I182 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2232), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I183 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .A(b_man[12]), .B(b_man[11]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I184 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060), .A(b_man[13]), .B(b_man[11]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I185 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3060), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I186 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947), .A(b_man[13]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I187 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I188 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3449), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3152), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3041));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I189 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I190 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3381), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I191 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I192 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3240), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I193 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I194 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I195 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3039), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2910), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2639));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I196 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I197 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3112), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I198 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2914), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I199 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I200 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2775), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2576), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3158));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I201 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3640), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2793));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I202 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2856), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2456), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2312));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I203 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3075), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3214), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3687));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I204 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3100), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I205 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .A(a_man[10]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I206 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I207 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .A(a_man[11]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I209 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2230), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I210 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3448));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I211 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I212 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3502), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I213 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8352));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I214 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I215 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2432), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I216 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I217 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2296), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I218 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I219 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2572), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I220 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3643), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3504), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2225));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I221 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3425), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3172), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2889));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I222 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I223 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2841), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I224 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I225 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2703), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I226 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712), .A(b_man[10]), .B(b_man[9]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I227 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I228 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I229 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267), .A(b_man[11]), .B(b_man[9]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I230 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2267), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2712));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I231 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258), .A(b_man[11]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I232 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I233 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2495), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2363), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2817));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I234 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3109), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3025), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3306));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I235 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2515), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3580), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2716));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I236 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3663), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2256), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2739));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2415), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I238 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3307), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I242 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3444), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I244 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2706), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2972), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3107));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I246 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3173), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I247 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3110), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I248 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I249 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2843), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2774), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2426));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I250 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2462), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2319), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3606));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I251 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2549), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3247), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2371));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I252 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3520), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2174), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2531));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I253 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3293), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I254 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .A(a_man[8]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I255 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .A(a_man[9]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I257 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I258 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2429), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I259 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3641));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I260 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I261 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2634), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I262 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I263 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2497), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2768), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I266 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2291), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2159), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2425));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I267 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3648), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3117), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2574));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I268 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2689), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3084), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3670));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I270 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2157), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3570), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I273 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3371), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3234), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3527));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I275 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3032), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I276 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2902), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I278 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2218), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I280 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3637), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I283 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2356), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I284 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3438), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3300), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3562));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I285 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2564), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2556));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2364), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I288 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779), .A(b_man[8]), .B(b_man[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I289 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I290 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I291 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033), .A(b_man[9]), .B(b_man[7]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I292 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3033), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2779));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I293 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564), .A(b_man[9]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I294 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I295 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2473), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3140));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3498), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3373), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I300 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I301 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I302 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3168), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3035), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2772));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I303 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I304 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3237), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I305 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3305), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I306 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I307 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2903), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2970), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3250));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I308 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3092), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3286), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2884));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I309 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3255), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3313), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2782));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I310 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2202), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2605), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3279));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I311 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2149), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2289), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3294));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I312 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2617), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I313 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2965), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2836), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I317 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I318 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3099), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I319 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2626), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2490), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2762));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I320 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I321 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2567), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I322 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I323 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2428), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2699), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I326 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2222), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3639), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2359));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I327 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2870), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3398));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I328 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2918), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2973), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2209));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I329 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3340), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2262), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2376));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I330 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2747), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3365), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3496));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I331 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I332 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .A(a_man[6]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I333 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I334 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .A(a_man[7]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I335 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I336 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2631), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I337 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2288));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I338 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2756), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3408), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2951));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I339 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2435), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2696), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3589));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I340 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2944), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2522), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2309));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2821), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844), .A(b_man[6]), .B(b_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I345 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242), .A(b_man[7]), .B(b_man[5]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2242), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2844));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332), .A(b_man[7]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I349 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I350 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3227), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I351 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I353 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I354 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I358 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I360 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2829), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2693), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2956));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I362 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8328));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I366 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I367 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I368 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I369 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I370 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I371 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2418), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2287), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2559));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I372 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I373 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I374 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3439), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2765), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I375 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3567), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2894), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I376 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2838), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3103), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3229));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I377 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2276), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2819), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2924));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I378 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3680), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2893), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3038));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I379 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3064), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3380), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2405));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I380 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .A(a_man[4]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I382 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .A(a_man[5]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I384 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I385 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2487));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2557), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I388 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2284), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3164), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I389 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2153), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3028), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I390 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2417), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3292), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I391 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3492), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3366), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3630));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I392 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3354), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2210), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3179));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I393 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3303), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2629), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I394 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3497), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2835), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I396 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2967), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3167), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2785));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I397 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3506), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3235), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2668));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I398 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3203), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2644), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2187));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I399 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3431), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3149));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I400 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3534), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2530), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2358));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I401 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3501), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3372), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2181));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2493), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906), .A(b_man[4]), .B(b_man[3]));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I406 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I407 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004), .A(b_man[5]), .B(b_man[3]));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3004), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2906));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I409 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645), .A(b_man[5]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I411 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2156), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3350), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2446));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I412 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I413 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3430), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I414 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2351), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2214), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2483), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I420 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3556), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3432), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3689));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I421 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3093), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2798), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3479));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I422 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3015), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2901), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3484));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I423 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3633), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I425 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I426 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3495), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I427 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I428 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I429 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3297), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3166), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2897));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I431 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3368), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I432 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2150), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I433 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I434 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3030), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3364), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2824));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I435 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3328), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3511), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2190));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I436 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2299), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2475), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2705));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I437 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3675), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2790), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3458));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I438 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2610), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3031), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3171));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I439 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3014), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I440 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I441 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2757), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I442 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I443 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2618), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .A(a_man[2]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I446 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .A(a_man[3]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3026), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I449 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2690));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I450 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2408), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2277), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2625));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I451 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3094), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I454 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2957), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I455 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I456 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3223), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I457 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2758), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2623), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2890));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I458 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8320));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I459 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I460 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2695), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I461 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I462 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2562), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I463 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I464 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2833), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I465 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2354), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2216), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2484));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I466 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3106), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3636), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2961));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I467 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2679), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2252), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2449));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I468 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2986), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3184), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2708));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I469 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3155), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3463), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3683));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I470 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2441), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2416), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3098));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I471 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2813), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3596), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2154));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I472 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2339), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I473 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968), .A(b_man[2]), .B(b_man[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I474 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211), .A(b_man[3]), .B(b_man[1]));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I477 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2211), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2968));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I478 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959), .A(b_man[3]));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I480 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3482), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I483 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3362), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I485 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3622), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I486 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3156), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3021), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3287));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I487 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3012), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2285), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3517));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I488 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I489 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2686), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I490 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I491 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2554), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I492 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I493 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2820), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I494 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2345), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2206), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2474));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I495 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I496 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2279), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I498 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2148), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2410), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I501 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3485), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3363), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3625));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I502 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3216), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2198), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2486));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I503 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2227), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2571), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3302));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I504 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2349), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I505 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .A(a_man[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I506 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I507 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I508 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3554), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3370));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I509 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I510 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I511 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I512 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3434), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I513 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3558), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I515 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2962), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3096), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3226));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I516 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2602), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2742), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2229));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I517 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3658), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2770), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3132));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I518 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3629), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2391), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3071));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I519 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2563), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3125), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3265));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I520 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3209), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I522 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3289), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I524 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3160), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I525 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3426), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I527 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2952), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2822), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3087));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I528 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I529 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2892), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I530 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2760), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I533 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3023), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I534 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2555), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2411), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2688));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I535 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2915), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3252));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I536 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I537 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3684), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I539 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3550), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I540 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I541 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I542 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I543 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3355), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3217), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3476));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I544 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I545 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2624), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I546 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3220), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I548 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2282), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2887), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2641));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I549 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2518), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2778), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3500));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I550 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2950), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2270), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I551 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2611), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2258), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2997));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I552 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3420), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2396), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2883));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I553 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3605), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3575), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2735));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I554 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2763), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3210), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3230));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I555 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2538), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I556 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .A(a_man[0]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I557 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I558 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I559 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272), .A(b_man[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I561 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .A(b_man[0]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I562 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
NAND2X2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I563 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I565 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3085), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2350));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807), .A(b_man[21]), .B(b_man[22]));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I567 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I568 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2807), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2400));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I569 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I570 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8295));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I571 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I573 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I575 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I576 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2479), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2616));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I577 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I578 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2476), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I579 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2348), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I581 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I582 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2613), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I583 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3686), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3551), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2272));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I584 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2724), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2183), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3602));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I585 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I586 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I587 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I588 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3478), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I590 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I592 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I593 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3282), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3151), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3419));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I594 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I595 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3219), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I596 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I597 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I598 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I599 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8336));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I600 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I601 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3358), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I602 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2886), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2754), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3016));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I603 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2691));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I604 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3627), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2954), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I605 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2207), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3089), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I606 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3024), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3291), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3428));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I607 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2666), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3199), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2306));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I608 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2550), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3423), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I609 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3488), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2825), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I610 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2203), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2748), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3162));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I611 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I612 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3150), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I613 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2882), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2199), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I614 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2751), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3618), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I615 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I616 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3013), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I617 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2545), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2403), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2680));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I618 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3086), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2814), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3353));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I619 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3555), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2553), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3027));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I620 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I621 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2178), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2677), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2431));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I622 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3367), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2353), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2789));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I623 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3427), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2891), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2528));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I624 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3192), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2579), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3585));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I625 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3078), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2661), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2746));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I626 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3443), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2424), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2346));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I627 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2964), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2685), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3274));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I628 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2170), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3242), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2876));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I629 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3414), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I630 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I631 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I632 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I633 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I634 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3079), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I635 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2877), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2743), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3228));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I636 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I637 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2546), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I638 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I639 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2406), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I640 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I641 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2683), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I642 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2201), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3620), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2341));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I643 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3316), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2496), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2828));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I644 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I645 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2816), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I646 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I647 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I648 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I649 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I650 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2946), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I651 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2470), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3005), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2606));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I652 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I653 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3688), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I654 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2799), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I655 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3553), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I656 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I657 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2274), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I658 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3361), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3221), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3480));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I659 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2638), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3034), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3076));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I660 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2338), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3211), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I661 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3538), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2379), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2570));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I662 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2864), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3402), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2322));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I663 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2234), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2837), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2268));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I664 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3611), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2316));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I665 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2831), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2909), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3389));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I666 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2734), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I667 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I668 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3284), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I669 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I670 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3153), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I671 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I672 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3422), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I673 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2949), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2818), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3080));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I674 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I675 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3678), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I676 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I677 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3542), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I678 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I679 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2264), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I680 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3348), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3213), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3472));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I681 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2333), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3347), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2290));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I682 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2468), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3346), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I683 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2452), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I684 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2888), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I685 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I686 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3019), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I687 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2548), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2684));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I688 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I689 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2537), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I690 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I691 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2397), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I692 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I693 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2673), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I694 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2192), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3612), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2330));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I695 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3205), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2815), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3584));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I696 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2698), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3676), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2158));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I697 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3222), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2810), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3097));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I698 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3249), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2859), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2489));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I699 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2803), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3549), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2482));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I700 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3604), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I701 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3530), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3057), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2525));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I702 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2692), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2205), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3473));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I703 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3521), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2971), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2457));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I704 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I705 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I706 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3276), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I707 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I708 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3146), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I709 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I710 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3413), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I711 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2941), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2811), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3070));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I712 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2872), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2247), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2551));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I713 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2975), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2297), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2471));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I714 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I715 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2472), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I716 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I717 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2343), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I718 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I719 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2609), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I720 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3681), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3545), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2266));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I721 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I722 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2879), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I723 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I724 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2745), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I725 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I726 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3008), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I727 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2539), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2399), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2675));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I728 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3323), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2794), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2809));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I729 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3375), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3009), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2360));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I730 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2465), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3454), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2585));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I731 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2633), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3617), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2152));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I732 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I733 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529), .A(b_man[19]), .B(b_man[20]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I734 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871), .A(b_man[21]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2529));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I735 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3660), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I736 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2204), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I737 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2871), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3424));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I738 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I739 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2736), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I740 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I741 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2600), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I742 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595), .A(b_man[17]), .B(b_man[18]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I743 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933), .A(b_man[19]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2595));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I744 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3329), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I745 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2987), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I746 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I747 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2933), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3615));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I748 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2392), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2259), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2878));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I749 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3533), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2385), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2395), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3609));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I750 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3384), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3204), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2980));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I751 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2648), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2386));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I752 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3083), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2401), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I753 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I754 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3215), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I755 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2749), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2880));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I756 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2764), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2303), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3315));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I757 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I758 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2334), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I759 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I760 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2194), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I761 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I762 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2463), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I763 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3535), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3416), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3672));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I764 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I765 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3474), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I766 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I767 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3351), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I768 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I769 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3613), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I770 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3147), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3010), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3278));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I771 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3236), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2221), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3563));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I772 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3459), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2443), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3677));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I773 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3119), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2953), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3624));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I774 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3590), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3145), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3281));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I775 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I776 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I777 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3072), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I778 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I779 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2942), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I780 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I781 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3206), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I782 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2738), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2603), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2873));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I783 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2420), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3357), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2532));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I784 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I785 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3468), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I786 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I787 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3342), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I788 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3603), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2450), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2993), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2659));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I789 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3137), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2999), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3271));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I790 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I791 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2541), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I792 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I793 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2812), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I794 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I795 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2678), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I796 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2196), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2467), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2335));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I797 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3487), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2340), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2791));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I798 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2905), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3441), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3599));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I799 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3066), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2674), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2612));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I800 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2241), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2213), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3335));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I801 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I802 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I803 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3673), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I804 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I805 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3537), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I806 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I807 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2261), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I808 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3345), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3207), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3470));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I809 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I810 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2533), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I811 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I812 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2393), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I813 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I814 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2667), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I815 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2189), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3607), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2323));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I816 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2654), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3661), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3541));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I817 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2653), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I818 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3280), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I819 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I820 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3417), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I821 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2943), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3074));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I822 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3514), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2540), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3295));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I823 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3544), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3042), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3018));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I824 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3128), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3654), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2504));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I825 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2534), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3288), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3433));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I826 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I827 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658), .A(b_man[15]), .B(b_man[16]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I828 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994), .A(b_man[17]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2658));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I829 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2308), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I830 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2604), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I831 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2994), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2263));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I832 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I833 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2804), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I834 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2628), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2458), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3187));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I835 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I836 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2874), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I837 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I838 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2740), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8298), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I839 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I840 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3003), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I841 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2535), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2394), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2669));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I842 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I843 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3273), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I844 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I845 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3141), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I846 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I847 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3410), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I848 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2937), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2806), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3065));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I849 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3304), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2773), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2253));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I850 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2254), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3159), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3330));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I851 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2566), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3102), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2622));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I852 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2730), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3508), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3056));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I853 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I854 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I855 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3528), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8358), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I856 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3665), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2519), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3583), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2860));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I857 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3513), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I858 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3471), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I859 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I860 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3608), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I861 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3143), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3275));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I862 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3200), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3336), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2200));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I863 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2310), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2912), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3464));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I864 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3212), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2936), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2682));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I865 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2164), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3632), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2271));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I866 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I867 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2966), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2286), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2575));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I868 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I869 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2731), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I870 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I871 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2596), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I872 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I873 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2865), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I874 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2387), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2255), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2523));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I875 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I876 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2328), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I877 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I878 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2191), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I879 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I880 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2460), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I881 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3532), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3411), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3667));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I882 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2687), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3218), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2512));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I883 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3579), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2427), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2988));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I884 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3073), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2278), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3040));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I885 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I886 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721), .A(b_man[13]), .B(b_man[14]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I887 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058), .A(b_man[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2721));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I888 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I889 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2808), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I890 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3058), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2461));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I891 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3338), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3421), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2771));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I892 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I893 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3465), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I894 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I895 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3339), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I896 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I897 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3597), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I898 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3133), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2996), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3267));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I899 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I900 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3067), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I901 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I902 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2939), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I903 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I904 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3201), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I905 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2733), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2598), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2869));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I906 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2260), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2805), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3022));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I907 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2347), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2885), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3244));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I908 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2172), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2597), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2737));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I909 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I910 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I911 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2184), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8359), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2352), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2923));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I912 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2853), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I913 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3669), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I914 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I915 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2257), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I916 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3341), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3466));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I917 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3403), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3450), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3277));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I918 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I919 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2526), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I920 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I921 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2390), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I922 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I923 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2662), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I924 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2185), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3600), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2318));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I925 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2581), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2995), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3522));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I926 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2459), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2547));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I927 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2832), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3638), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3392));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I928 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I929 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I930 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I931 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I932 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I933 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3524), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I934 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I935 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2947), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I936 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3331), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3193), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3460));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I937 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I938 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3268), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I939 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I940 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3135), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I941 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I942 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3406), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8325), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I943 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2932), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2802), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3062));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I944 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3113), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2492));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I945 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2929), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2646), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2248), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2981));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I946 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2800), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8342), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3659), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I947 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795), .A(b_man[11]), .B(b_man[12]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I948 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126), .A(b_man[13]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2795));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I949 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2511), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I950 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2998), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I951 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3126), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2664));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I952 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2592), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2453), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3369));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I953 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3399), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2719), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3668));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I954 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2398), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3552), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2485));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I955 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I956 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I957 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I958 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2725), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I959 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I960 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2594), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I961 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I962 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2861), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I963 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2383), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2249), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2520));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I964 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3029), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3429), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2235));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I965 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2374), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2236), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3169));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I966 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3523), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3142), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3614));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I967 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I968 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2171), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I969 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2321), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I970 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I971 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2455), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I972 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3525), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3662));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I973 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855), .A(b_man[9]), .B(b_man[10]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I974 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185), .A(b_man[11]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2855));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I975 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3391), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I976 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3195), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I977 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3185), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2863));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I978 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I979 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2989), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I980 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2311), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8343), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3258), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3048));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I981 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I982 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2179), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8334), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I983 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3047), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I984 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2521), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I985 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I986 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I987 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I988 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2180), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2314));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I989 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3515), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3400), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2382));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I990 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3002), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2652), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2608));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I991 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2155), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2407), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3557));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I992 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3644), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3052), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3194));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I993 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I994 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I995 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I996 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3462), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I997 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3334), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2655), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I998 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I999 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3593), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1000 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3129), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2991), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3261));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1001 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3619), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2466), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2491));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1002 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2839), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3088), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3311));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1003 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1004 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1005 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2927), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1006 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1007 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2796), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1008 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1009 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3053), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1010 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2589), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2448), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2718));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1011 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3061), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2671), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2752));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1012 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3225), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3674), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2753));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1013 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1014 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1015 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916), .A(b_man[7]), .B(b_man[8]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1016 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251), .A(b_man[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2916));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1017 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2713), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1018 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3401), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1019 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3251), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3054));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1020 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1021 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3655), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1022 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1023 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3519), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1024 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1025 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2243), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1026 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3324), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3188), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3457));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1027 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3592), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3121), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2245));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1028 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3202), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2265), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3344));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1029 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1030 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2368), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1031 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2720), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1032 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1033 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2858), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1034 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2378), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2517));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1035 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2375), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8335), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3564), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3114));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1036 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3174), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3586), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2788));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1037 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2727), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3263), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2868));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1038 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1039 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1040 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1041 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3122), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1042 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1043 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2984), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1044 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978), .A(b_man[5]), .B(b_man[6]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1045 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317), .A(b_man[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2978));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1046 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3578), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1047 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3588), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1048 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3317), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3253));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1049 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2786), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2649), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3037));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1050 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3319), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3456), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3001));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1051 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1052 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1053 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1054 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2305), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1055 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1056 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2173), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1057 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2440), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8327), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2332), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3175));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1058 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3510), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3396), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3650));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1059 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2499), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2846), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2977));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1060 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1061 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3243), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1062 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2920), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1063 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1064 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3051), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1065 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2584), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2715));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1066 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3231), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2700), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3260));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1067 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1068 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045), .A(b_man[3]), .B(b_man[4]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1069 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385), .A(b_man[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3045));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1070 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2911), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1071 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2237), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1072 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3385), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3452));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1073 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1074 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3183), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1075 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3436), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2850), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2899));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1076 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1077 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1078 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2507), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8310), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2645), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2302));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1079 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1080 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2370), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1081 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2573), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1082 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3116), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1083 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1084 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3246), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1085 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2781), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2913));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1086 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2166), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3582), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2759));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1087 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1088 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1089 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1090 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111), .A(b_man[1]), .B(b_man[2]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1091 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446), .A(b_man[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3111));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1092 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2228), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1093 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2437), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
ADDHX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1094 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3446), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3647));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1095 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1096 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2577), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8302), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2959), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2620));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1097 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1098 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1099 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1100 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3312), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
OAI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1101 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2636), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2357), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3272), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2935));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1102 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1103 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1104 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2231), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3290));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1105 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1106 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2769), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2423));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1107 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3626), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2412));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1108 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1109 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3095), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2215));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1110 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1111 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3574), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3241));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1112 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2561), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3569));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1113 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1114 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2362), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3377));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1115 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1116 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2650), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2307));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1117 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2161), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3649));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1118 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2439), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2588));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1119 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505));
AOI31X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1120 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176), .A2(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3270));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1121 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2926), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3531));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1122 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1123 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3539), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3208));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1124 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2327), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2948));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1125 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3283), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2355));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1126 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1127 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2414), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3628));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1128 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2694), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2433));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1129 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2780), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2317));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1130 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244));
OAI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1131 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2621), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2281));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1132 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2663), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2744));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1133 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3082), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3165));
AO21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1134 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1135 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3264), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2928));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1136 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2513));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1137 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2854), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3415));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1138 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1139 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1140 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2193), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2960));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1141 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2842), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527));
OAI31X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1142 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3148), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160), .A2(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3091));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1143 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3296), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2849));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1144 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2578));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1145 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3182), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3409));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1146 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3397));
OAI2BB2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1147 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2188), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2558));
OAI2BB2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1148 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2896), .B1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2922));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1149 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3259), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2404));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1150 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2741));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1151 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2750), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3309));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1152 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3547));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1153 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3642), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3139));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1154 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2827));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1155 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3467), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3163));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1156 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3144), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2934), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3254), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3635));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1157 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2908), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3491), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2508));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1158 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151), .A0N(N11566), .A1N(N11564), .B0(N11830));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1159 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2168), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2852), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3540));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1160 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393), .A0N(N11560), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151), .B0(N11822));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1161 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2985), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2337), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3437));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1162 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197), .A0N(N11554), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393), .B0(N11814));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1163 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2250), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2220), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2384));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1164 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239), .A0N(N11548), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197), .B0(N11806));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1165 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3069), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2729), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3477));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1166 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412), .A0N(N11542), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239), .B0(N11798));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1167 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2336), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2269), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2293));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1168 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701), .A0N(N11536), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412), .B0(N11790));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1169 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3154), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2637), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2862));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1170 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670), .A0N(N11530), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701), .B0(N11782));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1171 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2413), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3196), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3616));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1172 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310), .A0N(N11524), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670), .B0(N11774));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1173 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3233), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2402), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2630));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1174 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081), .A0N(N11518), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310), .B0(N11766));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1175 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2501), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2969), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3049));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1176 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516), .A0N(N11512), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081), .B0(N11758));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1177 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3320), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2992));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1178 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104), .A0N(N11506), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516), .B0(N11750));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1179 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2591), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3332), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3418));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1180 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349), .A0N(N11500), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104), .B0(N11742));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1181 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3407), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2195), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2826));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1182 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723), .A0N(N11177), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349), .B0(N11734));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1183 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2672), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3161), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2421));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1184 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776), .A0N(N11171), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723), .B0(N11726));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1185 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3475), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3044), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2767));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1186 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493), .A0N(N11165), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776), .B0(N11718));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1187 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2755), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3386), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3656));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1188 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356), .A0N(N11159), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493), .B0(N11710));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1189 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3561), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2447), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3601));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1190 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331), .A0N(N11153), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356), .B0(N11702));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1191 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2840), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2389));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1192 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526), .A0N(N11147), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331), .B0(N11694));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1193 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3645), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3352), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2875));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1194 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315), .A0N(N11141), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526), .B0(N11686));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1195 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2917), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2275), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3679));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1196 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326), .A0N(N11135), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315), .B0(N11678));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1197 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2320), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2963));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1198 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2938), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3134));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1199 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3178), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2614), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2761));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1200 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3326), .B(N11675));
BUFX2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1201 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47]));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1202 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1203 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1204 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2315), .B(N11135));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1205 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1206 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3356), .B(N11153));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1207 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2331), .B(N11147));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1208 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1209 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3493), .B(N11159));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1210 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[43]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1211 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1212 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3526), .B(N11141));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1213 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[46]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1214 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[44]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[45]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1215 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1216 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5370));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1217 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3393), .B(N11554));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1218 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2197), .B(N11548));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1219 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8368));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1220 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1221 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2151), .B(N11560));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1222 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[29]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1223 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1224 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27]), .A(N11564), .B(N11566));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1225 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[28]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1226 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26]), .A(N11570), .B(N11572));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1227 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[27]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1228 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1229 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5405), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1230 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[25]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2494), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2251));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1231 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26]), .A(N11241), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[26]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1232 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2409), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3131));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1233 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]), .A(N11239), .B(N11241), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1234 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1235 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[23]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3007), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2451));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1236 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24]), .A(N10847), .B(N11239), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1237 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1238 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5411), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]));
NAND2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1239 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5378), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1240 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3516), .B(N11506));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1241 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3104), .B(N11500));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1242 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1243 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3081), .B(N11512));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1244 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[37]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1245 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1246 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3310), .B(N11518));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1247 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[36]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1248 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2670), .B(N11524));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1249 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[35]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1250 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1251 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5345), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1252 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2701), .B(N11530));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1253 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[34]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1254 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3412), .B(N11536));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1255 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[33]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1256 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1257 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3239), .B(N11542));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1258 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[32]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1259 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[30]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[31]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1260 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1261 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5390), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1262 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5412), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1263 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8402));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1264 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2776), .B(N11165));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1265 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[42]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1266 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2723), .B(N11171));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1267 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[41]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1268 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1269 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3349), .B(N11177));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1270 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[40]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1271 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[38]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[39]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1272 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1273 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5408), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1274 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5337), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1275 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[47]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8411));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1276 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2728), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3327));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1277 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23]), .A(N10845), .B(N10847), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1278 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1279 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1280 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23), .A(a_sign), .B(b_sign));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1281 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N445), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1282 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1283 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1284 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N446), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1285 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2640), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2976));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1286 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2834), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2660));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1287 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1288 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3666));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1289 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10]), .A(N11364), .B(N11366), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1290 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1291 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3560), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1292 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2244), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2590));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1293 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3006), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3610));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1294 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1295 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3077));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1296 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14]), .A(N11385), .B(N11387), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1297 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3651), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2514), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3318));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1298 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2438), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2787));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1299 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3360), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3138));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1300 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3123), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3455));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1301 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2478), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2601));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1302 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12]), .A(N11406), .B(N11408), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1303 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3262), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2445), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2925));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1304 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3594), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2381));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1305 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2895), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2543));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1306 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1307 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3548));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1308 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16]), .A(N11343), .B(N11345), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1309 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[10]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[14]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[12]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[16]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1310 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3435), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2217));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1311 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2560), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2898));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1312 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2326), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3308));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1313 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2]), .A(N11350), .B(N11352), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1314 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3036), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3376));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1315 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3170), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3248));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1316 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2162), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2498));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1317 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2582), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2717));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1318 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6]), .A(N11359), .B(N11373), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1319 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3232), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3568));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1320 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2607), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2777));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1321 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2361), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2702));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1322 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2208), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2233));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1323 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4]), .A(N11392), .B(N11357), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1324 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1325 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2177));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1326 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3176), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3337), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2845));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1327 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3505), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2298));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1328 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2147), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3191));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1329 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8]), .A(N11401), .B(N11378), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1330 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[6]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[4]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[8]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1331 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5528), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5538));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1332 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5]), .A(N11357), .B(N11359), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1333 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9]), .A(N11378), .B(N11364), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1334 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7]), .A(N11373), .B(N11401), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1335 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11]), .A(N11366), .B(N11406), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1336 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[5]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[9]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[7]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[11]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1337 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3]), .A(N11352), .B(N11392), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1338 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3124), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2651));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1339 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22]), .A(N11449), .B(N10845), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1340 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[22]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1341 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3388), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2851));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1342 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2643), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3512));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1343 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20]), .A(N11454), .B(N11447), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1344 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3063));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1345 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2726));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1346 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3621), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3285));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1347 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3405), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2186));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1348 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3020));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1349 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2160), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3565), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3374));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1350 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2527), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2867));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1351 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N3224), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2481));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1352 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18]), .A(N11468), .B(N11470), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1353 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[20]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[18]));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1354 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[0]), .A(b_man[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2292));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1355 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376), .B(N11475));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1356 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1]), .A(N11475), .B(N11350), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8376));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1357 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21]), .A(N11447), .B(N11449), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8373));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1358 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19]), .A(N11470), .B(N11454), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1359 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17]), .A(N11345), .B(N11468), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1360 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[19]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[17]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1361 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15]), .A(N11387), .B(N11343), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1362 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13]), .A(N11408), .B(N11385), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5224));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1363 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[15]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[13]));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1364 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5536), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5547));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1365 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[1]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[21]), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5545));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1366 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5530), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5540), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5558));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1367 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5554), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5532));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1368 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5552), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5543));
NOR3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1369 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
OA21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1370 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[24]), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34), .B0(N10872));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1371 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447), .A(N10827), .B(N10829), .C(N10831), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N444));
OAI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1372 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450), .A0(N10829), .A1(N10831), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__34));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1373 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[23]), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N447), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N450));
AOI21X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1374 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[24]), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__24[47]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1375 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0]), .A(N10694), .B(N10696), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1376 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631), .A(b_exp[0]), .B(a_exp[0]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1377 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]), .A(b_exp[1]), .B(a_exp[1]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5631));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1378 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1379 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]), .A(b_exp[2]), .B(a_exp[2]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5624));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1380 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1381 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[2]), .A(N10703), .B(N10705), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1382 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]), .A(b_exp[3]), .B(a_exp[3]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5643));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1383 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5697));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1384 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1385 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]), .A(b_exp[4]), .B(a_exp[4]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5655));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1386 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1387 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[4]), .A(N10712), .B(N10714), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1388 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1389 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]), .A(b_exp[5]), .B(a_exp[5]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5637));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1390 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5681), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1391 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[5]), .A(N10721), .B(N10723), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1392 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812), .A(N10621), .B(N10623), .C(N10625), .D(N10627));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1393 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]), .A(b_exp[6]), .B(a_exp[6]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5652));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1394 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[4]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[5]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5701));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1395 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1396 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627), .A(a_exp[7]));
ADDFX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1397 (.CO(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647), .S(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5627), .B(b_exp[7]), .CI(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5632));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1398 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5699), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1399 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[7]), .A(N10739), .B(N10741), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1400 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5682), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[3]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1401 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[3]), .A(N10757), .B(N10759), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
AND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1402 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1403 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8]), .A(a_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1404 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1405 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[8]), .A(N10774), .B(N10776), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1406 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[1]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1407 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[1]), .A(N10766), .B(N10768), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1408 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813), .A(N10616), .B(N11432));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1409 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5700), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[6]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1410 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[6]), .A(N10748), .B(N10750), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1411 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5691));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1412 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]), .A(a_exp[7]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5647));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1413 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__31[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5690), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1414 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[9]), .A(N10730), .B(N10732), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__38));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1415 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801), .A(N11425), .B(N10643));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1416 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5813), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5801));
NOR3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1417 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808), .A(N10630), .B(N10632), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5815));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1418 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__20), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__13));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1419 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__21), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__14));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1420 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830), .A(N10637), .B(N10639), .C(N10490), .D(N10643));
OAI2BB1X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1421 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823), .A0N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5812), .A1N(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5808), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5830));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1422 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768), .A(N11432), .B(N11425));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1423 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763), .A(N10630), .B(N10632));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1424 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775), .A(N10625), .B(N10623));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1425 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772), .A(N10621), .B(N10627));
NOR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1426 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5768), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5763), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5775), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5772));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1427 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417), .A(N10616), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N461));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1428 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8417), .B(N10643));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1429 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5823), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__51));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1430 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1431 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .A(N10438), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1432 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10262));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1433 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1434 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5366), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]));
AND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1435 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028), .A(N10412), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6695 (.Y(N13001), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6028));
INVX2 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6696 (.Y(N13002), .A(N13001));
NOR2BX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1436 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887), .B(N10412));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1437 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951), .A0(N10146), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10152));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1438 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6014), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1439 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380), .A(N10464), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
INVX1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6697 (.Y(N13003), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8380));
INVX3 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I6698 (.Y(N13004), .A(N13003));
NOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1440 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .A(N10490), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1441 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852), .A(rm[0]), .B(rm[1]));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1442 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7), .A(rm[2]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5852));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1443 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__7), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__6));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1444 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5860), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5500), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__5));
OR4X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1445 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1446 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[8]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[7]));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1447 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__30[9]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N442));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1448 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5914), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1449 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043), .A0(N9948), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1450 (.Y(x[21]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6048), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5951), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6043));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1451 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10257));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1452 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1453 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5400), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[44]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1454 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061), .A0(N10137), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10143));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1455 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069), .A0(N9939), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1456 (.Y(x[20]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5965), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6061), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6069));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1457 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10252));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1458 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1459 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5341), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[43]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1460 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977), .A0(N10128), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10134));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1461 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091), .A0(N9930), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1462 (.Y(x[19]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6075), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5977), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6091));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1463 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10247));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1464 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1465 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5369), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[42]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1466 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084), .A0(N10119), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10125));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1467 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117), .A0(N9921), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1468 (.Y(x[18]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5990), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6084), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6117));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1469 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10242));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1470 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5422), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1471 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5404), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[41]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1472 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002), .A0(N10110), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10116));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1473 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948), .A0(N9912), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1474 (.Y(x[17]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6098), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6002), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5948));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1475 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10237));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1476 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1477 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5344), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[40]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1478 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109), .A0(N10101), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10107));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1479 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973), .A0(N9903), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1480 (.Y(x[16]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6016), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6109), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5973));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1481 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10232));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1482 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[39]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1483 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027), .A0(N10092), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10098));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1484 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999), .A0(N9894), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1485 (.Y(x[15]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5931), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6027), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5999));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1486 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10227));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1487 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1488 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5419), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1489 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5394), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[38]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1490 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941), .A0(N10083), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10089));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1491 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024), .A0(N9885), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1492 (.Y(x[14]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6038), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5941), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6024));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1493 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10222));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1494 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5353), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1495 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5359), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[37]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1496 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051), .A0(N10074), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10080));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1497 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047), .A0(N9876), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1498 (.Y(x[13]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5955), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6051), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6047));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1499 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10217));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1500 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1501 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5351), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[36]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1502 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967), .A0(N10065), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10071));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1503 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073), .A0(N9867), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1504 (.Y(x[12]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6063), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5967), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6073));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1505 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10212));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1506 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5365));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1507 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5333), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[35]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1508 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077), .A0(N10056), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10062));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1509 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096), .A0(N9858), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1510 (.Y(x[11]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5980), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6077), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6096));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1511 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10207));
NOR3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1512 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1513 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5363), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[34]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1514 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992), .A0(N10047), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10053));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1515 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930), .A0(N9849), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1516 (.Y(x[10]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6086), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5992), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5930));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1517 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10202));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1518 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5403), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1519 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5385), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[33]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1520 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100), .A0(N10038), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10044));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1521 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953), .A0(N9840), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1522 (.Y(x[9]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6005), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6100), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5953));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1523 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10197));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1524 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1525 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5361), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[32]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1526 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018), .A0(N10029), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10035));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1527 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978), .A0(N9831), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1528 (.Y(x[8]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6112), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6018), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5978));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1529 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10192));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1530 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5373), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[31]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1531 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933), .A0(N10020), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10026));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1532 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004), .A0(N9822), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1533 (.Y(x[7]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6032), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5933), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6004));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1534 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10187));
NAND3BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1535 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1536 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5406), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[30]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1537 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040), .A0(N10011), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10017));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1538 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030), .A0(N9813), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1539 (.Y(x[6]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5943), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6040), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6030));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1540 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10182));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1541 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5416), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1542 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5346), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[29]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1543 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957), .A0(N10002), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N10008));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1544 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053), .A0(N9804), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1545 (.Y(x[5]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6055), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5957), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6053));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1546 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10177));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1547 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1548 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5375), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[28]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1549 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066), .A0(N9993), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N9999));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1550 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079), .A0(N9795), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1551 (.Y(x[4]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5970), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6066), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6079));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1552 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10172));
XOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1553 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5387), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[27]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1554 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982), .A0(N9984), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N9990));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1555 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102), .A0(N9786), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1556 (.Y(x[3]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6080), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5982), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6102));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1557 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10167));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1558 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1559 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5338), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[26]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1560 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088), .A0(N9975), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N9981));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1561 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934), .A0(N9777), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1562 (.Y(x[2]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5996), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6088), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5934));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1563 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10162));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1564 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[0]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[25]));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1565 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008), .A0(N9966), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N9972));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1566 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959), .A0(N9768), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1567 (.Y(x[1]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6104), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6008), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5959));
NAND2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1568 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8382), .B(N10157));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1569 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114), .A0(N9957), .A1(N13002), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5987), .B1(N9963));
AOI22XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1570 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984), .A0(N9759), .A1(N13004), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N8378), .B1(N13000));
NAND3XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1571 (.Y(x[0]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6020), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N6114), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5984));
NAND4BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1572 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336), .AN(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5371), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[45]), .C(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5392), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5384));
XNOR2X1 float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1573 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5336), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1574 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5923), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__25[46]), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[22]), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__44));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1575 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5925), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__47));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1576 (.Y(x[22]), .A(N9514), .B(N9512), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__49));
NOR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1577 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__28), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__32));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1578 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__27), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26));
OR2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1579 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5874), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1580 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5887));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1581 (.Y(x[30]), .A(N10630), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1582 (.Y(x[29]), .A(N11425), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1583 (.Y(x[28]), .A(N10627), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1584 (.Y(x[27]), .A(N10625), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1585 (.Y(x[26]), .A(N10632), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1586 (.Y(x[25]), .A(N10623), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1587 (.Y(x[24]), .A(N11432), .B(N9467), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
INVXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1588 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5870), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__48[0]));
AOI21XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1589 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5893), .A0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__42), .A1(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N469), .B0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N470));
MXI2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1590 (.Y(x[23]), .A(N9507), .B(N9505), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N5884));
NAND2BXL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1591 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135), .AN(b_sign), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__22));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1592 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2135), .B(a_sign), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__15));
MX2XL float_div_cynw_cm_float_mul_ieee_E8_M23_4_I1593 (.Y(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31]), .A(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__23), .B(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_N2140), .S0(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__26));
EDFFHQX1 x_reg_L0_31__I1625 (.Q(N4032), .D(float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[31]), .E(bdw_enable), .CK(aclk));
EDFFHQX1 x_reg_L1_31__I1657 (.Q(x[31]), .D(N4032), .E(bdw_enable), .CK(aclk));
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[0] = x[0];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[1] = x[1];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[2] = x[2];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[3] = x[3];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[4] = x[4];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[5] = x[5];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[6] = x[6];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[7] = x[7];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[8] = x[8];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[9] = x[9];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[10] = x[10];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[11] = x[11];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[12] = x[12];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[13] = x[13];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[14] = x[14];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[15] = x[15];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[16] = x[16];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[17] = x[17];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[18] = x[18];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[19] = x[19];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[20] = x[20];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[21] = x[21];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[22] = x[22];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[23] = x[23];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[24] = x[24];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[25] = x[25];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[26] = x[26];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[27] = x[27];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[28] = x[28];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[29] = x[29];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_x[30] = x[30];
assign float_div_cynw_cm_float_mul_ieee_E8_M23_2_inst_inst_cellmath__45[23] = 1'B0;
endmodule

/* CADENCE  vbnwTArcoh4= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



