/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:11:00 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_2_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__9,
	inst_cellmath__17;
wire [8:0] inst_cellmath__19;
wire [7:0] inst_cellmath__20;
wire [8:0] inst_cellmath__22;
wire  inst_cellmath__28,
	inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__33,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42;
wire [15:0] inst_cellmath__48;
wire [18:0] inst_cellmath__51;
wire [24:0] inst_cellmath__60;
wire [39:0] inst_cellmath__62__W0, inst_cellmath__62__W1,
	inst_cellmath__63__W0, inst_cellmath__63__W1;
wire [39:0] inst_cellmath__64;
wire  inst_cellmath__67;
wire N446,N447,N448,N449,N450,N451,N452 
	,N453,N454,N455,N456,N457,N458,N477,N478 
	,N479,N480,N481,N482,N483,N484,N485,N486 
	,N487,N488,N489,N490,N491,N492,N493,N494 
	,N495,N496,N497,N498,N499,N500,N501;
cynw_cm_float_rcp_inst_cellmath__9_0_bdw1412651405_bdw cynw_cm_float_rcp_I0 (.inst_cellmath__9_0_out0(inst_cellmath__9), .inst_cellmath__9_0_in0({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_rcp_inst_cellmath__15__5__bdw1412651405_bdw cynw_cm_float_rcp_I1 (.inst_cellmath__15__5__out0(inst_cellmath__19[0]), .inst_cellmath__15__5__in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16], a_man[15], a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_rcp_inst_cellmath__29_0_bdw1412651405_bdw cynw_cm_float_rcp_I2 (.inst_cellmath__29_0_out0(inst_cellmath__29), .inst_cellmath__29_0_in0(inst_cellmath__9), .inst_cellmath__29_0_in1(inst_cellmath__19[0]));
cynw_cm_float_rcp_inst_cellmath__37_0_bdw1412651405_bdw cynw_cm_float_rcp_I3 (.inst_cellmath__37_0_out0(x[31]), .inst_cellmath__37_0_in0(inst_cellmath__29), .inst_cellmath__37_0_in1(a_sign));
cynw_cm_float_rcp_inst_cellmath__28_0_bdw1412651405_bdw cynw_cm_float_rcp_I4 (.inst_cellmath__28_0_out0(inst_cellmath__28), .inst_cellmath__28_0_in0(inst_cellmath__9), .inst_cellmath__28_0_in1(inst_cellmath__19[0]));
INVXL cynw_cm_float_rcp_I5 (.Y(inst_cellmath__20[0]), .A(a_exp[0]));
INVXL cynw_cm_float_rcp_I6 (.Y(inst_cellmath__20[1]), .A(a_exp[1]));
INVXL cynw_cm_float_rcp_I7 (.Y(inst_cellmath__20[2]), .A(a_exp[2]));
INVXL cynw_cm_float_rcp_I8 (.Y(inst_cellmath__20[3]), .A(a_exp[3]));
INVXL cynw_cm_float_rcp_I9 (.Y(inst_cellmath__20[4]), .A(a_exp[4]));
INVXL cynw_cm_float_rcp_I10 (.Y(inst_cellmath__20[5]), .A(a_exp[5]));
INVXL cynw_cm_float_rcp_I11 (.Y(inst_cellmath__20[6]), .A(a_exp[6]));
INVXL cynw_cm_float_rcp_I12 (.Y(inst_cellmath__20[7]), .A(a_exp[7]));
cynw_cm_float_rcp_inst_cellmath__22_0_bdw1412651405_bdw cynw_cm_float_rcp_I13 (.inst_cellmath__22_0_out0({inst_cellmath__22[8], inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}), .inst_cellmath__22_0_in0({inst_cellmath__20[7], inst_cellmath__20[6], inst_cellmath__20[5], inst_cellmath__20[4], inst_cellmath__20[3], inst_cellmath__20[2], inst_cellmath__20[1], inst_cellmath__20[0]}), .inst_cellmath__22_0_in1(inst_cellmath__19[0]));
cynw_cm_float_rcp_inst_cellmath__17__6__bdw1412651405_bdw cynw_cm_float_rcp_I14 (.inst_cellmath__17__6__out0({N446}), .inst_cellmath__17__6__in0({inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}));
cynw_cm_float_rcp_inst_cellmath__17_0_bdw1412651405_bdw cynw_cm_float_rcp_I15 (.inst_cellmath__17_0_out0(inst_cellmath__17), .inst_cellmath__17_0_in0({inst_cellmath__22[8]}), .inst_cellmath__17_0_in1({N446}));
cynw_cm_float_rcp_inst_cellmath__30_0_bdw1412651405_bdw cynw_cm_float_rcp_I16 (.inst_cellmath__30_0_out0(inst_cellmath__30), .inst_cellmath__30_0_in0(inst_cellmath__9), .inst_cellmath__30_0_in1(inst_cellmath__17));
cynw_cm_float_rcp_inst_cellmath__33__7__bdw1412651405_bdw cynw_cm_float_rcp_I17 (.inst_cellmath__33__7__out0({N447}), .inst_cellmath__33__7__in0(inst_cellmath__30), .inst_cellmath__33__7__in1(inst_cellmath__28));
cynw_cm_float_rcp_inst_cellmath__33_0_bdw1412651405_bdw cynw_cm_float_rcp_I18 (.inst_cellmath__33_0_out0(inst_cellmath__33), .inst_cellmath__33_0_in0({N447}), .inst_cellmath__33_0_in1(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__34_0_bdw1412651405_bdw cynw_cm_float_rcp_I19 (.inst_cellmath__34_0_out0(inst_cellmath__34), .inst_cellmath__34_0_in0(inst_cellmath__29), .inst_cellmath__34_0_in1({a_exp[7], a_exp[6], a_exp[5], a_exp[4], a_exp[3], a_exp[2], a_exp[1], a_exp[0]}));
cynw_cm_float_rcp_inst_cellmath__42__9__bdw1412651405_bdw cynw_cm_float_rcp_I20 (.inst_cellmath__42__9__out0(inst_cellmath__42), .inst_cellmath__42__9__in0(inst_cellmath__34), .inst_cellmath__42__9__in1(inst_cellmath__33), .inst_cellmath__42__9__in2(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__38_0_bdw1412651405_bdw cynw_cm_float_rcp_I21 (.inst_cellmath__38_0_out0(inst_cellmath__38), .inst_cellmath__38_0_in0(inst_cellmath__34), .inst_cellmath__38_0_in1(inst_cellmath__29));
cynw_cm_float_rcp_inst_cellmath__43_0_bdw1412651405_bdw cynw_cm_float_rcp_I22 (.inst_cellmath__43_0_out0({x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23]}), .inst_cellmath__43_0_in0(inst_cellmath__42), .inst_cellmath__43_0_in1(inst_cellmath__38), .inst_cellmath__43_0_in2({inst_cellmath__22[7], inst_cellmath__22[6], inst_cellmath__22[5], inst_cellmath__22[4], inst_cellmath__22[3], inst_cellmath__22[2], inst_cellmath__22[1], inst_cellmath__22[0]}));
cynw_cm_float_rcp_inst_cellmath__67__11__bdw1412651405_bdw cynw_cm_float_rcp_I23 (.inst_cellmath__67__11__out0({N448}), .inst_cellmath__67__11__in0(inst_cellmath__34), .inst_cellmath__67__11__in1(inst_cellmath__33), .inst_cellmath__67__11__in2(inst_cellmath__29), .inst_cellmath__67__11__in3(inst_cellmath__19[0]));
INVXL cynw_cm_float_rcp_I24 (.Y(inst_cellmath__67), .A(N448));
INVXL cynw_cm_float_rcp_I25 (.Y(inst_cellmath__48[15]), .A(a_man[15]));
cynw_cm_float_rcp_inst_cellmath__60_0_bdw1412651405_bdw cynw_cm_float_rcp_I26 (.inst_cellmath__60_0_out0({inst_cellmath__60[24], inst_cellmath__60[23], inst_cellmath__60[22], inst_cellmath__60[21], inst_cellmath__60[20], inst_cellmath__60[19], inst_cellmath__60[18], inst_cellmath__60[17], inst_cellmath__60[16], inst_cellmath__60[15], inst_cellmath__60[14], inst_cellmath__60[13], inst_cellmath__60[12], inst_cellmath__60[11], inst_cellmath__60[10], inst_cellmath__60[9], inst_cellmath__60[8], inst_cellmath__60[7], inst_cellmath__60[6], inst_cellmath__60[5], inst_cellmath__60[4], inst_cellmath__60[3], inst_cellmath__60[2], inst_cellmath__60[1], inst_cellmath__60[0]}), .inst_cellmath__60_0_in0(inst_cellmath__48[15]), .inst_cellmath__60_0_in1({a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3]}));
cynw_cm_float_rcp_inst_noninc_a_cellmath__55_2WWMM_bdw1412651405_bdw cynw_cm_float_rcp_I27 (.inst_noninc_a_cellmath__55_2WWMM_out0({N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, inst_cellmath__51[17], inst_cellmath__51[16], inst_cellmath__51[15], inst_cellmath__51[14], inst_cellmath__51[13], inst_cellmath__51[12], inst_cellmath__51[11], inst_cellmath__51[10], inst_cellmath__51[9], inst_cellmath__51[8], inst_cellmath__51[7], inst_cellmath__51[6], inst_cellmath__51[5], inst_cellmath__51[4], inst_cellmath__51[3], inst_cellmath__51[2], inst_cellmath__51[1], inst_cellmath__51[0], N458, N457, N456, N455, N454, N453, N452, N451, N450, N449}), .inst_noninc_a_cellmath__55_2WWMM_in0({a_man[22], a_man[21], a_man[20], a_man[19], a_man[18], a_man[17], a_man[16]}));
cynw_cm_float_rcp_inst_cellmath__62_0_bdw1412651405_bdw cynw_cm_float_rcp_I28 (.inst_cellmath__62_0_out0({inst_cellmath__62__W1[39], inst_cellmath__62__W1[38], inst_cellmath__62__W1[37], inst_cellmath__62__W1[36], inst_cellmath__62__W1[35], inst_cellmath__62__W1[34], inst_cellmath__62__W1[33], inst_cellmath__62__W1[32], inst_cellmath__62__W1[31], inst_cellmath__62__W1[30], inst_cellmath__62__W1[29], inst_cellmath__62__W1[28], inst_cellmath__62__W1[27], inst_cellmath__62__W1[26], inst_cellmath__62__W1[25], inst_cellmath__62__W1[24], inst_cellmath__62__W1[23], inst_cellmath__62__W1[22], inst_cellmath__62__W1[21], inst_cellmath__62__W1[20], inst_cellmath__62__W1[19], inst_cellmath__62__W1[18], inst_cellmath__62__W1[17], inst_cellmath__62__W1[16], inst_cellmath__62__W1[15], inst_cellmath__62__W1[14], inst_cellmath__62__W1[13], inst_cellmath__62__W1[12], inst_cellmath__62__W1[11], inst_cellmath__62__W1[10], inst_cellmath__62__W1[9], inst_cellmath__62__W1[8], inst_cellmath__62__W1[7], inst_cellmath__62__W1[6], inst_cellmath__62__W1[5], inst_cellmath__62__W1[4], inst_cellmath__62__W1[3], inst_cellmath__62__W1[2], inst_cellmath__62__W1[1], inst_cellmath__62__W1[0]}), .inst_cellmath__62_0_out1({inst_cellmath__62__W0[39], inst_cellmath__62__W0[38], inst_cellmath__62__W0[37], inst_cellmath__62__W0[36], inst_cellmath__62__W0[35], inst_cellmath__62__W0[34], inst_cellmath__62__W0[33], inst_cellmath__62__W0[32], inst_cellmath__62__W0[31], inst_cellmath__62__W0[30], inst_cellmath__62__W0[29], inst_cellmath__62__W0[28], inst_cellmath__62__W0[27], inst_cellmath__62__W0[26], inst_cellmath__62__W0[25], inst_cellmath__62__W0[24], inst_cellmath__62__W0[23], inst_cellmath__62__W0[22], inst_cellmath__62__W0[21], inst_cellmath__62__W0[20], inst_cellmath__62__W0[19], inst_cellmath__62__W0[18], inst_cellmath__62__W0[17], inst_cellmath__62__W0[16], inst_cellmath__62__W0[15], inst_cellmath__62__W0[14], inst_cellmath__62__W0[13], inst_cellmath__62__W0[12], inst_cellmath__62__W0[11], inst_cellmath__62__W0[10], inst_cellmath__62__W0[9], inst_cellmath__62__W0[8], inst_cellmath__62__W0[7], inst_cellmath__62__W0[6], inst_cellmath__62__W0[5], inst_cellmath__62__W0[4], inst_cellmath__62__W0[3], inst_cellmath__62__W0[2], inst_cellmath__62__W0[1], inst_cellmath__62__W0[0]}), .inst_cellmath__62_0_in0({N458, N457, N456, N455, N454, N453, N452, N451, N450, N449}), .inst_cellmath__62_0_in1({inst_cellmath__60[24], inst_cellmath__60[23], inst_cellmath__60[22], inst_cellmath__60[21], inst_cellmath__60[20], inst_cellmath__60[19], inst_cellmath__60[18], inst_cellmath__60[17], inst_cellmath__60[16], inst_cellmath__60[15], inst_cellmath__60[14], inst_cellmath__60[13]}));
cynw_cm_float_rcp_inst_cellmath__63_0_bdw1412651405_bdw cynw_cm_float_rcp_I29 (.inst_cellmath__63_0_out0({inst_cellmath__63__W1[39], inst_cellmath__63__W1[38], inst_cellmath__63__W1[37], inst_cellmath__63__W1[36], inst_cellmath__63__W1[35], inst_cellmath__63__W1[34], inst_cellmath__63__W1[33], inst_cellmath__63__W1[32], inst_cellmath__63__W1[31], inst_cellmath__63__W1[30], inst_cellmath__63__W1[29], inst_cellmath__63__W1[28], inst_cellmath__63__W1[27], inst_cellmath__63__W1[26], inst_cellmath__63__W1[25], inst_cellmath__63__W1[24], inst_cellmath__63__W1[23], inst_cellmath__63__W1[22], inst_cellmath__63__W1[21], inst_cellmath__63__W1[20], inst_cellmath__63__W1[19], inst_cellmath__63__W1[18], inst_cellmath__63__W1[17], inst_cellmath__63__W1[16], inst_cellmath__63__W1[15], inst_cellmath__63__W1[14], inst_cellmath__63__W1[13], inst_cellmath__63__W1[12], inst_cellmath__63__W1[11], inst_cellmath__63__W1[10], inst_cellmath__63__W1[9], inst_cellmath__63__W1[8], inst_cellmath__63__W1[7], inst_cellmath__63__W1[6], inst_cellmath__63__W1[5], inst_cellmath__63__W1[4], inst_cellmath__63__W1[3], inst_cellmath__63__W1[2], inst_cellmath__63__W1[1], inst_cellmath__63__W1[0]}), .inst_cellmath__63_0_out1({inst_cellmath__63__W0[39], inst_cellmath__63__W0[38], inst_cellmath__63__W0[37], inst_cellmath__63__W0[36], inst_cellmath__63__W0[35], inst_cellmath__63__W0[34], inst_cellmath__63__W0[33], inst_cellmath__63__W0[32], inst_cellmath__63__W0[31], inst_cellmath__63__W0[30], inst_cellmath__63__W0[29], inst_cellmath__63__W0[28], inst_cellmath__63__W0[27], inst_cellmath__63__W0[26], inst_cellmath__63__W0[25], inst_cellmath__63__W0[24], inst_cellmath__63__W0[23], inst_cellmath__63__W0[22], inst_cellmath__63__W0[21], inst_cellmath__63__W0[20], inst_cellmath__63__W0[19], inst_cellmath__63__W0[18], inst_cellmath__63__W0[17], inst_cellmath__63__W0[16], inst_cellmath__63__W0[15], inst_cellmath__63__W0[14], inst_cellmath__63__W0[13], inst_cellmath__63__W0[12], inst_cellmath__63__W0[11], inst_cellmath__63__W0[10], inst_cellmath__63__W0[9], inst_cellmath__63__W0[8], inst_cellmath__63__W0[7], inst_cellmath__63__W0[6], inst_cellmath__63__W0[5], inst_cellmath__63__W0[4], inst_cellmath__63__W0[3], inst_cellmath__63__W0[2], inst_cellmath__63__W0[1], inst_cellmath__63__W0[0]}), .inst_cellmath__63_0_in0({inst_cellmath__51[17], inst_cellmath__51[16], inst_cellmath__51[15], inst_cellmath__51[14], inst_cellmath__51[13], inst_cellmath__51[12], inst_cellmath__51[11], inst_cellmath__51[10], inst_cellmath__51[9], inst_cellmath__51[8], inst_cellmath__51[7], inst_cellmath__51[6], inst_cellmath__51[5], inst_cellmath__51[4], inst_cellmath__51[3], inst_cellmath__51[2], inst_cellmath__51[1], inst_cellmath__51[0]}), .inst_cellmath__63_0_in1(inst_cellmath__48[15]), .inst_cellmath__63_0_in2({a_man[14], a_man[13], a_man[12], a_man[11], a_man[10], a_man[9], a_man[8], a_man[7], a_man[6], a_man[5], a_man[4], a_man[3], a_man[2], a_man[1], a_man[0]}));
cynw_cm_float_rcp_inst_cellmath__64_0_bdw1412651405_bdw cynw_cm_float_rcp_I30 (.inst_cellmath__64_0_out0({inst_cellmath__64[39], inst_cellmath__64[38], inst_cellmath__64[37], inst_cellmath__64[36], inst_cellmath__64[35], inst_cellmath__64[34], inst_cellmath__64[33], inst_cellmath__64[32], inst_cellmath__64[31], inst_cellmath__64[30], inst_cellmath__64[29], inst_cellmath__64[28], inst_cellmath__64[27], inst_cellmath__64[26], inst_cellmath__64[25], inst_cellmath__64[24], inst_cellmath__64[23], inst_cellmath__64[22], inst_cellmath__64[21], inst_cellmath__64[20], inst_cellmath__64[19], inst_cellmath__64[18], inst_cellmath__64[17], inst_cellmath__64[16], inst_cellmath__64[15], inst_cellmath__64[14], inst_cellmath__64[13], inst_cellmath__64[12], inst_cellmath__64[11], inst_cellmath__64[10], inst_cellmath__64[9], inst_cellmath__64[8], inst_cellmath__64[7], inst_cellmath__64[6], inst_cellmath__64[5], inst_cellmath__64[4], inst_cellmath__64[3], inst_cellmath__64[2], inst_cellmath__64[1], inst_cellmath__64[0]}), .inst_cellmath__64_0_in0({N501, N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477}), .inst_cellmath__64_0_in1({inst_cellmath__63__W1[39], inst_cellmath__63__W1[38], inst_cellmath__63__W1[37], inst_cellmath__63__W1[36], inst_cellmath__63__W1[35], inst_cellmath__63__W1[34], inst_cellmath__63__W1[33], inst_cellmath__63__W1[32], inst_cellmath__63__W1[31], inst_cellmath__63__W1[30], inst_cellmath__63__W1[29], inst_cellmath__63__W1[28], inst_cellmath__63__W1[27], inst_cellmath__63__W1[26], inst_cellmath__63__W1[25], inst_cellmath__63__W1[24], inst_cellmath__63__W1[23], inst_cellmath__63__W1[22], inst_cellmath__63__W1[21], inst_cellmath__63__W1[20], inst_cellmath__63__W1[19], inst_cellmath__63__W1[18], inst_cellmath__63__W1[17], inst_cellmath__63__W1[16], inst_cellmath__63__W1[15], inst_cellmath__63__W1[14], inst_cellmath__63__W1[13], inst_cellmath__63__W1[12], inst_cellmath__63__W1[11], inst_cellmath__63__W1[10], inst_cellmath__63__W1[9], inst_cellmath__63__W1[8], inst_cellmath__63__W1[7], inst_cellmath__63__W1[6], inst_cellmath__63__W1[5], inst_cellmath__63__W1[4], inst_cellmath__63__W1[3], inst_cellmath__63__W1[2], inst_cellmath__63__W1[1], inst_cellmath__63__W1[0]}), .inst_cellmath__64_0_in2({inst_cellmath__63__W0[39], inst_cellmath__63__W0[38], inst_cellmath__63__W0[37], inst_cellmath__63__W0[36], inst_cellmath__63__W0[35], inst_cellmath__63__W0[34], inst_cellmath__63__W0[33], inst_cellmath__63__W0[32], inst_cellmath__63__W0[31], inst_cellmath__63__W0[30], inst_cellmath__63__W0[29], inst_cellmath__63__W0[28], inst_cellmath__63__W0[27], inst_cellmath__63__W0[26], inst_cellmath__63__W0[25], inst_cellmath__63__W0[24], inst_cellmath__63__W0[23], inst_cellmath__63__W0[22], inst_cellmath__63__W0[21], inst_cellmath__63__W0[20], inst_cellmath__63__W0[19], inst_cellmath__63__W0[18], inst_cellmath__63__W0[17], inst_cellmath__63__W0[16], inst_cellmath__63__W0[15], inst_cellmath__63__W0[14], inst_cellmath__63__W0[13], inst_cellmath__63__W0[12], inst_cellmath__63__W0[11], inst_cellmath__63__W0[10], inst_cellmath__63__W0[9], inst_cellmath__63__W0[8], inst_cellmath__63__W0[7], inst_cellmath__63__W0[6], inst_cellmath__63__W0[5], inst_cellmath__63__W0[4], inst_cellmath__63__W0[3], inst_cellmath__63__W0[2], inst_cellmath__63__W0[1], inst_cellmath__63__W0[0]}), .inst_cellmath__64_0_in3({inst_cellmath__62__W1[39], inst_cellmath__62__W1[38], inst_cellmath__62__W1[37], inst_cellmath__62__W1[36], inst_cellmath__62__W1[35], inst_cellmath__62__W1[34], inst_cellmath__62__W1[33], inst_cellmath__62__W1[32], inst_cellmath__62__W1[31], inst_cellmath__62__W1[30], inst_cellmath__62__W1[29], inst_cellmath__62__W1[28], inst_cellmath__62__W1[27], inst_cellmath__62__W1[26], inst_cellmath__62__W1[25], inst_cellmath__62__W1[24], inst_cellmath__62__W1[23], inst_cellmath__62__W1[22], inst_cellmath__62__W1[21], inst_cellmath__62__W1[20], inst_cellmath__62__W1[19], inst_cellmath__62__W1[18], inst_cellmath__62__W1[17], inst_cellmath__62__W1[16], inst_cellmath__62__W1[15], inst_cellmath__62__W1[14], inst_cellmath__62__W1[13], inst_cellmath__62__W1[12], inst_cellmath__62__W1[11], inst_cellmath__62__W1[10], inst_cellmath__62__W1[9], inst_cellmath__62__W1[8], inst_cellmath__62__W1[7], inst_cellmath__62__W1[6], inst_cellmath__62__W1[5], inst_cellmath__62__W1[4], inst_cellmath__62__W1[3], inst_cellmath__62__W1[2], inst_cellmath__62__W1[1], inst_cellmath__62__W1[0]}), .inst_cellmath__64_0_in4({inst_cellmath__62__W0[39], inst_cellmath__62__W0[38], inst_cellmath__62__W0[37], inst_cellmath__62__W0[36], inst_cellmath__62__W0[35], inst_cellmath__62__W0[34], inst_cellmath__62__W0[33], inst_cellmath__62__W0[32], inst_cellmath__62__W0[31], inst_cellmath__62__W0[30], inst_cellmath__62__W0[29], inst_cellmath__62__W0[28], inst_cellmath__62__W0[27], inst_cellmath__62__W0[26], inst_cellmath__62__W0[25], inst_cellmath__62__W0[24], inst_cellmath__62__W0[23], inst_cellmath__62__W0[22], inst_cellmath__62__W0[21], inst_cellmath__62__W0[20], inst_cellmath__62__W0[19], inst_cellmath__62__W0[18], inst_cellmath__62__W0[17], inst_cellmath__62__W0[16], inst_cellmath__62__W0[15], inst_cellmath__62__W0[14], inst_cellmath__62__W0[13], inst_cellmath__62__W0[12], inst_cellmath__62__W0[11], inst_cellmath__62__W0[10], inst_cellmath__62__W0[9], inst_cellmath__62__W0[8], inst_cellmath__62__W0[7], inst_cellmath__62__W0[6], inst_cellmath__62__W0[5], inst_cellmath__62__W0[4], inst_cellmath__62__W0[3], inst_cellmath__62__W0[2], inst_cellmath__62__W0[1], inst_cellmath__62__W0[0]}));
cynw_cm_float_rcp_inst_cellmath__68_0_bdw1412651405_bdw cynw_cm_float_rcp_I31 (.inst_cellmath__68_0_out0({x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .inst_cellmath__68_0_in0(inst_cellmath__67), .inst_cellmath__68_0_in1({inst_cellmath__64[39], inst_cellmath__64[38], inst_cellmath__64[37], inst_cellmath__64[36], inst_cellmath__64[35], inst_cellmath__64[34], inst_cellmath__64[33], inst_cellmath__64[32], inst_cellmath__64[31], inst_cellmath__64[30], inst_cellmath__64[29], inst_cellmath__64[28], inst_cellmath__64[27], inst_cellmath__64[26], inst_cellmath__64[25], inst_cellmath__64[24], inst_cellmath__64[23], inst_cellmath__64[22], inst_cellmath__64[21], inst_cellmath__64[20], inst_cellmath__64[19], inst_cellmath__64[18], inst_cellmath__64[17]}), .inst_cellmath__68_0_in2(inst_cellmath__29));
assign inst_cellmath__19[1] = 1'B1;
assign inst_cellmath__19[2] = 1'B1;
assign inst_cellmath__19[3] = 1'B1;
assign inst_cellmath__19[4] = 1'B1;
assign inst_cellmath__19[5] = 1'B1;
assign inst_cellmath__19[6] = 1'B1;
assign inst_cellmath__19[7] = 1'B1;
assign inst_cellmath__19[8] = 1'B1;
assign inst_cellmath__48[0] = a_man[0];
assign inst_cellmath__48[1] = a_man[1];
assign inst_cellmath__48[2] = a_man[2];
assign inst_cellmath__48[3] = a_man[3];
assign inst_cellmath__48[4] = a_man[4];
assign inst_cellmath__48[5] = a_man[5];
assign inst_cellmath__48[6] = a_man[6];
assign inst_cellmath__48[7] = a_man[7];
assign inst_cellmath__48[8] = a_man[8];
assign inst_cellmath__48[9] = a_man[9];
assign inst_cellmath__48[10] = a_man[10];
assign inst_cellmath__48[11] = a_man[11];
assign inst_cellmath__48[12] = a_man[12];
assign inst_cellmath__48[13] = a_man[13];
assign inst_cellmath__48[14] = a_man[14];
assign inst_cellmath__51[18] = 1'B1;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_cellmath__9_0_bdw1412651405_bdw (
	inst_cellmath__9_0_out0,
	inst_cellmath__9_0_in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__9_0_out0;
input [7:0] inst_cellmath__9_0_in0;
wire N11,N12,N13,N14,N15,N16;
NAND2XL inst_cellmath__9_0_I0 (.Y(N11), .A(inst_cellmath__9_0_in0[7]), .B(inst_cellmath__9_0_in0[0]));
NAND2XL inst_cellmath__9_0_I1 (.Y(N12), .A(inst_cellmath__9_0_in0[6]), .B(inst_cellmath__9_0_in0[5]));
NAND2XL inst_cellmath__9_0_I2 (.Y(N13), .A(inst_cellmath__9_0_in0[4]), .B(inst_cellmath__9_0_in0[3]));
NAND2XL inst_cellmath__9_0_I3 (.Y(N14), .A(inst_cellmath__9_0_in0[2]), .B(inst_cellmath__9_0_in0[1]));
NOR2XL inst_cellmath__9_0_I4 (.Y(N15), .A(N11), .B(N12));
NOR2XL inst_cellmath__9_0_I5 (.Y(N16), .A(N13), .B(N14));
AND2XL inst_cellmath__9_0_I6 (.Y(inst_cellmath__9_0_out0), .A(N15), .B(N16));
endmodule

module cynw_cm_float_rcp_inst_cellmath__15__5__bdw1412651405_bdw (
	inst_cellmath__15__5__out0,
	inst_cellmath__15__5__in0
	); /* architecture "gate_level" */ 
output  inst_cellmath__15__5__out0;
input [22:0] inst_cellmath__15__5__in0;
wire N27,N28,N29,N30,N31,N32,N33 
	,N34,N35,N36,N39,N40,N41,N44,N45 
	,N47,N48;
NOR2XL inst_cellmath__15__5__I1 (.Y(N27), .A(inst_cellmath__15__5__in0[22]), .B(inst_cellmath__15__5__in0[21]));
NOR2XL inst_cellmath__15__5__I2 (.Y(N28), .A(inst_cellmath__15__5__in0[20]), .B(inst_cellmath__15__5__in0[19]));
NOR2XL inst_cellmath__15__5__I3 (.Y(N29), .A(inst_cellmath__15__5__in0[18]), .B(inst_cellmath__15__5__in0[17]));
NOR2XL inst_cellmath__15__5__I4 (.Y(N30), .A(inst_cellmath__15__5__in0[16]), .B(inst_cellmath__15__5__in0[15]));
NOR2XL inst_cellmath__15__5__I5 (.Y(N31), .A(inst_cellmath__15__5__in0[14]), .B(inst_cellmath__15__5__in0[13]));
NOR2XL inst_cellmath__15__5__I6 (.Y(N32), .A(inst_cellmath__15__5__in0[12]), .B(inst_cellmath__15__5__in0[11]));
NOR2XL inst_cellmath__15__5__I7 (.Y(N33), .A(inst_cellmath__15__5__in0[10]), .B(inst_cellmath__15__5__in0[9]));
NOR2XL inst_cellmath__15__5__I8 (.Y(N34), .A(inst_cellmath__15__5__in0[8]), .B(inst_cellmath__15__5__in0[7]));
NOR2XL inst_cellmath__15__5__I9 (.Y(N35), .A(inst_cellmath__15__5__in0[6]), .B(inst_cellmath__15__5__in0[5]));
NOR2XL inst_cellmath__15__5__I10 (.Y(N36), .A(inst_cellmath__15__5__in0[4]), .B(inst_cellmath__15__5__in0[3]));
NAND2XL inst_cellmath__15__5__I13 (.Y(N39), .A(N27), .B(N28));
NAND2XL inst_cellmath__15__5__I14 (.Y(N40), .A(N29), .B(N30));
NAND2XL inst_cellmath__15__5__I15 (.Y(N41), .A(N31), .B(N32));
NOR4X1 inst_cellmath__15__5__I25 (.Y(N44), .A(inst_cellmath__15__5__in0[0]), .B(inst_cellmath__15__5__in0[1]), .C(inst_cellmath__15__5__in0[2]), .D(N39));
NOR2XL inst_cellmath__15__5__I19 (.Y(N45), .A(N40), .B(N41));
NAND4XL inst_cellmath__15__5__I27 (.Y(N48), .A(N33), .B(N35), .C(N34), .D(N36));
NAND2XL inst_cellmath__15__5__I21 (.Y(N47), .A(N44), .B(N45));
NOR2XL inst_cellmath__15__5__I23 (.Y(inst_cellmath__15__5__out0), .A(N48), .B(N47));
endmodule

module cynw_cm_float_rcp_inst_cellmath__29_0_bdw1412651405_bdw (
	inst_cellmath__29_0_out0,
	inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__29_0_out0;
input  inst_cellmath__29_0_in0,
	inst_cellmath__29_0_in1;
NOR2BX1 inst_cellmath__29_0_I2 (.Y(inst_cellmath__29_0_out0), .AN(inst_cellmath__29_0_in0), .B(inst_cellmath__29_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__37_0_bdw1412651405_bdw (
	inst_cellmath__37_0_out0,
	inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__37_0_out0;
input  inst_cellmath__37_0_in0,
	inst_cellmath__37_0_in1;
NOR2BX1 inst_cellmath__37_0_I2 (.Y(inst_cellmath__37_0_out0), .AN(inst_cellmath__37_0_in1), .B(inst_cellmath__37_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__28_0_bdw1412651405_bdw (
	inst_cellmath__28_0_out0,
	inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__28_0_out0;
input  inst_cellmath__28_0_in0,
	inst_cellmath__28_0_in1;
AND2XL inst_cellmath__28_0_I0 (.Y(inst_cellmath__28_0_out0), .A(inst_cellmath__28_0_in0), .B(inst_cellmath__28_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__22_0_bdw1412651405_bdw (
	inst_cellmath__22_0_out0,
	inst_cellmath__22_0_in0,
	inst_cellmath__22_0_in1
	); /* architecture "gate_level" */ 
output [8:0] inst_cellmath__22_0_out0;
input [7:0] inst_cellmath__22_0_in0;
input  inst_cellmath__22_0_in1;
wire N64,N68,N72,N76,N80,N84,N88 
	;
ADDHX1 inst_cellmath__22_0_I19 (.CO(N64), .S(inst_cellmath__22_0_out0[0]), .A(inst_cellmath__22_0_in0[0]), .B(inst_cellmath__22_0_in1));
XNOR2X1 hap1_A_I28 (.Y(inst_cellmath__22_0_out0[1]), .A(inst_cellmath__22_0_in0[1]), .B(N64));
OR2XL hap1_A_I29 (.Y(N68), .A(inst_cellmath__22_0_in0[1]), .B(N64));
XNOR2X1 hap1_A_I30 (.Y(inst_cellmath__22_0_out0[2]), .A(inst_cellmath__22_0_in0[2]), .B(N68));
OR2XL hap1_A_I31 (.Y(N72), .A(inst_cellmath__22_0_in0[2]), .B(N68));
XNOR2X1 hap1_A_I32 (.Y(inst_cellmath__22_0_out0[3]), .A(inst_cellmath__22_0_in0[3]), .B(N72));
OR2XL hap1_A_I33 (.Y(N76), .A(inst_cellmath__22_0_in0[3]), .B(N72));
XNOR2X1 hap1_A_I34 (.Y(inst_cellmath__22_0_out0[4]), .A(inst_cellmath__22_0_in0[4]), .B(N76));
OR2XL hap1_A_I35 (.Y(N80), .A(inst_cellmath__22_0_in0[4]), .B(N76));
XNOR2X1 hap1_A_I36 (.Y(inst_cellmath__22_0_out0[5]), .A(inst_cellmath__22_0_in0[5]), .B(N80));
OR2XL hap1_A_I37 (.Y(N84), .A(inst_cellmath__22_0_in0[5]), .B(N80));
XNOR2X1 hap1_A_I38 (.Y(inst_cellmath__22_0_out0[6]), .A(inst_cellmath__22_0_in0[6]), .B(N84));
OR2XL hap1_A_I39 (.Y(N88), .A(inst_cellmath__22_0_in0[6]), .B(N84));
XNOR2X1 hap1_A_I40 (.Y(inst_cellmath__22_0_out0[7]), .A(inst_cellmath__22_0_in0[7]), .B(N88));
NOR2XL hap1_A_I41 (.Y(inst_cellmath__22_0_out0[8]), .A(inst_cellmath__22_0_in0[7]), .B(N88));
endmodule

module cynw_cm_float_rcp_inst_cellmath__17__6__bdw1412651405_bdw (
	inst_cellmath__17__6__out0,
	inst_cellmath__17__6__in0
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__17__6__out0;
input [7:0] inst_cellmath__17__6__in0;
wire N17,N19,N20;
NOR3XL inst_cellmath__17__6__I14 (.Y(N20), .A(inst_cellmath__17__6__in0[2]), .B(inst_cellmath__17__6__in0[3]), .C(inst_cellmath__17__6__in0[5]));
NOR2XL inst_cellmath__17__6__I6 (.Y(N17), .A(inst_cellmath__17__6__in0[6]), .B(inst_cellmath__17__6__in0[7]));
NOR4BX1 inst_cellmath__17__6__I15 (.Y(N19), .AN(N17), .B(inst_cellmath__17__6__in0[0]), .C(inst_cellmath__17__6__in0[4]), .D(inst_cellmath__17__6__in0[1]));
NAND2X6 inst_cellmath__17__6__I10 (.Y(inst_cellmath__17__6__out0[0]), .A(N20), .B(N19));
endmodule

module cynw_cm_float_rcp_inst_cellmath__17_0_bdw1412651405_bdw (
	inst_cellmath__17_0_out0,
	inst_cellmath__17_0_in0,
	inst_cellmath__17_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__17_0_out0;
input [8:8] inst_cellmath__17_0_in0;
input [0:0] inst_cellmath__17_0_in1;
NAND2BXL inst_cellmath__17_0_I2 (.Y(inst_cellmath__17_0_out0), .AN(inst_cellmath__17_0_in0[8]), .B(inst_cellmath__17_0_in1[0]));
endmodule

module cynw_cm_float_rcp_inst_cellmath__30_0_bdw1412651405_bdw (
	inst_cellmath__30_0_out0,
	inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__30_0_out0;
input  inst_cellmath__30_0_in0,
	inst_cellmath__30_0_in1;
NOR2BX1 inst_cellmath__30_0_I3 (.Y(inst_cellmath__30_0_out0), .AN(inst_cellmath__30_0_in1), .B(inst_cellmath__30_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__33__7__bdw1412651405_bdw (
	inst_cellmath__33__7__out0,
	inst_cellmath__33__7__in0,
	inst_cellmath__33__7__in1
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__33__7__out0;
input  inst_cellmath__33__7__in0,
	inst_cellmath__33__7__in1;
OR2XL inst_cellmath__33__7__I0 (.Y(inst_cellmath__33__7__out0[0]), .A(inst_cellmath__33__7__in1), .B(inst_cellmath__33__7__in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__33_0_bdw1412651405_bdw (
	inst_cellmath__33_0_out0,
	inst_cellmath__33_0_in0,
	inst_cellmath__33_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__33_0_out0;
input [0:0] inst_cellmath__33_0_in0;
input  inst_cellmath__33_0_in1;
NOR2BX1 inst_cellmath__33_0_I3 (.Y(inst_cellmath__33_0_out0), .AN(inst_cellmath__33_0_in0[0]), .B(inst_cellmath__33_0_in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__34_0_bdw1412651405_bdw (
	inst_cellmath__34_0_out0,
	inst_cellmath__34_0_in0,
	inst_cellmath__34_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__34_0_out0;
input  inst_cellmath__34_0_in0;
input [7:0] inst_cellmath__34_0_in1;
wire N12,N13,N14,N15,N19;
NOR2XL inst_cellmath__34_0_I0 (.Y(N12), .A(inst_cellmath__34_0_in1[0]), .B(inst_cellmath__34_0_in1[1]));
NOR2XL inst_cellmath__34_0_I1 (.Y(N13), .A(inst_cellmath__34_0_in1[7]), .B(inst_cellmath__34_0_in1[6]));
NOR2XL inst_cellmath__34_0_I2 (.Y(N14), .A(inst_cellmath__34_0_in1[5]), .B(inst_cellmath__34_0_in1[4]));
NOR2XL inst_cellmath__34_0_I3 (.Y(N15), .A(inst_cellmath__34_0_in1[3]), .B(inst_cellmath__34_0_in1[2]));
NAND4XL inst_cellmath__34_0_I10 (.Y(N19), .A(N12), .B(N14), .C(N13), .D(N15));
NOR2XL inst_cellmath__34_0_I8 (.Y(inst_cellmath__34_0_out0), .A(N19), .B(inst_cellmath__34_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__42__9__bdw1412651405_bdw (
	inst_cellmath__42__9__out0,
	inst_cellmath__42__9__in0,
	inst_cellmath__42__9__in1,
	inst_cellmath__42__9__in2
	); /* architecture "gate_level" */ 
output  inst_cellmath__42__9__out0;
input  inst_cellmath__42__9__in0,
	inst_cellmath__42__9__in1,
	inst_cellmath__42__9__in2;
NOR3XL inst_cellmath__42__9__I3 (.Y(inst_cellmath__42__9__out0), .A(inst_cellmath__42__9__in2), .B(inst_cellmath__42__9__in0), .C(inst_cellmath__42__9__in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__38_0_bdw1412651405_bdw (
	inst_cellmath__38_0_out0,
	inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1
	); /* architecture "gate_level" */ 
output  inst_cellmath__38_0_out0;
input  inst_cellmath__38_0_in0,
	inst_cellmath__38_0_in1;
OR2XL inst_cellmath__38_0_I0 (.Y(inst_cellmath__38_0_out0), .A(inst_cellmath__38_0_in1), .B(inst_cellmath__38_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__43_0_bdw1412651405_bdw (
	inst_cellmath__43_0_out0,
	inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1,
	inst_cellmath__43_0_in2
	); /* architecture "gate_level" */ 
output [7:0] inst_cellmath__43_0_out0;
input  inst_cellmath__43_0_in0,
	inst_cellmath__43_0_in1;
input [7:0] inst_cellmath__43_0_in2;
MX2XL inst_cellmath__43_0_I16 (.Y(inst_cellmath__43_0_out0[0]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[0]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I17 (.Y(inst_cellmath__43_0_out0[1]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[1]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I18 (.Y(inst_cellmath__43_0_out0[2]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[2]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I19 (.Y(inst_cellmath__43_0_out0[3]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[3]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I20 (.Y(inst_cellmath__43_0_out0[4]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[4]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I21 (.Y(inst_cellmath__43_0_out0[5]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[5]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I22 (.Y(inst_cellmath__43_0_out0[6]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[6]), .S0(inst_cellmath__43_0_in0));
MX2XL inst_cellmath__43_0_I23 (.Y(inst_cellmath__43_0_out0[7]), .A(inst_cellmath__43_0_in1), .B(inst_cellmath__43_0_in2[7]), .S0(inst_cellmath__43_0_in0));
endmodule

module cynw_cm_float_rcp_inst_cellmath__67__11__bdw1412651405_bdw (
	inst_cellmath__67__11__out0,
	inst_cellmath__67__11__in0,
	inst_cellmath__67__11__in1,
	inst_cellmath__67__11__in2,
	inst_cellmath__67__11__in3
	); /* architecture "gate_level" */ 
output [0:0] inst_cellmath__67__11__out0;
input  inst_cellmath__67__11__in0,
	inst_cellmath__67__11__in1,
	inst_cellmath__67__11__in2,
	inst_cellmath__67__11__in3;
OR4X1 inst_cellmath__67__11__I7 (.Y(inst_cellmath__67__11__out0[0]), .A(inst_cellmath__67__11__in3), .B(inst_cellmath__67__11__in2), .C(inst_cellmath__67__11__in0), .D(inst_cellmath__67__11__in1));
endmodule

module cynw_cm_float_rcp_inst_cellmath__60_0_bdw1412651405_bdw (
	inst_cellmath__60_0_out0,
	inst_cellmath__60_0_in0,
	inst_cellmath__60_0_in1
	); /* architecture "gate_level" */ 
output [24:0] inst_cellmath__60_0_out0;
input  inst_cellmath__60_0_in0;
input [14:3] inst_cellmath__60_0_in1;
wire N80,N84,N86,N88,N90,N92,N94 
	,N96,N98,N100,N118,N120,N122,N124,N126 
	,N128,N130,N132,N134,N136,N150,N154,N156 
	,N158,N160,N162,N164,N166,N168,N170,N184 
	,N188,N190,N192,N194,N196,N198,N200,N202 
	,N216,N220,N222,N224,N226,N228,N230,N232 
	,N246,N250,N252,N254,N256,N258,N260,N274 
	,N278,N280,N282,N284,N286,N300,N304,N306 
	,N308,N310,N324,N328,N330,N332,N346,N350 
	,N352,N366,N370,N384,N404,N405,N406,N407 
	,N408,N409,N410,N411,N412,N413,N414,N415 
	,N416,N417,N418,N419,N420,N421,N422,N423 
	,N424,N425,N426,N427,N428,N429,N430,N431 
	,N432,N433,N434,N435,N436,N437,N438,N439 
	,N440,N441,N442,N443,N444,N445,N446,N447 
	,N448,N449,N450,N451,N452,N453,N454,N455 
	,N456,N457,N458,N459,N460,N461,N462,N463 
	,N464,N465,N466,N469,N470,N471,N472,N473 
	,N474,N475,N476,N477,N478,N479,N480,N481 
	,N482,N483,N484,N485,N486,N487,N488,N489 
	,N490,N491,N492,N493,N494,N495,N496,N497 
	,N498,N499,N500,N501,N502,N503,N504,N505 
	,N506,N507,N508,N509,N510,N511,N512,N513 
	,N514,N515,N516,N517,N518,N519,N520,N521 
	,N522,N523,N524,N525,N526,N527,N528,N529 
	,N530,N531,N532,N533,N534,N535,N536,N537 
	,N538,N541,N551,N559,N571,N583,N611,N614 
	,N617,N620,N623,N632,N634,N635,N636,N637 
	,N638,N639,N640,N641,N642,N643,N644,N645 
	,N646,N647,N648,N649,N650,N651,N652,N653 
	,N654,N655,N656,N657,N658,N659,N660,N661 
	,N662,N663,N665,N668,N674,N682,N692,N704 
	,N718,N734,N752,N772,N794,N818,N844,N872 
	,N902,N934,N1170,N1171,N1172,N1183,N1184,N1190 
	,N1191,N1192,N1193,N1194,N1195,N1196,N1201,N1203 
	,N1204,N1210,N1211,N1221,N1222;
INVXL inst_cellmath__60_0_I761 (.Y(N1170), .A(inst_cellmath__60_0_in1[4]));
INVXL inst_cellmath__60_0_I762 (.Y(N1171), .A(inst_cellmath__60_0_in1[5]));
INVXL inst_cellmath__60_0_I763 (.Y(N1172), .A(inst_cellmath__60_0_in1[6]));
INVXL inst_cellmath__60_0_I774 (.Y(N1183), .A(inst_cellmath__60_0_in1[7]));
INVXL inst_cellmath__60_0_I775 (.Y(N1184), .A(inst_cellmath__60_0_in1[8]));
INVXL inst_cellmath__60_0_I781 (.Y(N1190), .A(inst_cellmath__60_0_in1[9]));
INVXL inst_cellmath__60_0_I782 (.Y(N1191), .A(inst_cellmath__60_0_in1[10]));
INVXL inst_cellmath__60_0_I783 (.Y(N1192), .A(inst_cellmath__60_0_in1[11]));
INVXL inst_cellmath__60_0_I784 (.Y(N1193), .A(inst_cellmath__60_0_in1[12]));
INVXL inst_cellmath__60_0_I785 (.Y(N1194), .A(inst_cellmath__60_0_in1[13]));
INVXL inst_cellmath__60_0_I786 (.Y(N1195), .A(inst_cellmath__60_0_in1[14]));
INVXL inst_cellmath__60_0_I787 (.Y(N1196), .A(inst_cellmath__60_0_in0));
INVXL inst_cellmath__60_0_I792 (.Y(N1201), .A(inst_cellmath__60_0_in1[3]));
OR2XL inst_cellmath__60_0_I1366 (.Y(N80), .A(N1201), .B(N1170));
NOR2XL inst_cellmath__60_0_I20 (.Y(N528), .A(N1201), .B(N1171));
NOR2XL inst_cellmath__60_0_I21 (.Y(N84), .A(N1201), .B(N1172));
NOR2XL inst_cellmath__60_0_I22 (.Y(N86), .A(N1201), .B(N1183));
NOR2XL inst_cellmath__60_0_I23 (.Y(N88), .A(N1201), .B(N1184));
NOR2XL inst_cellmath__60_0_I24 (.Y(N90), .A(N1201), .B(N1190));
NOR2XL inst_cellmath__60_0_I25 (.Y(N92), .A(N1201), .B(N1191));
NOR2XL inst_cellmath__60_0_I26 (.Y(N94), .A(N1201), .B(N1192));
NOR2XL inst_cellmath__60_0_I27 (.Y(N96), .A(N1201), .B(N1193));
NOR2XL inst_cellmath__60_0_I28 (.Y(N98), .A(N1201), .B(N1194));
NOR2XL inst_cellmath__60_0_I29 (.Y(N100), .A(N1201), .B(N1195));
OR2XL inst_cellmath__60_0_I30 (.Y(N404), .A(N1201), .B(N1196));
NOR2XL inst_cellmath__60_0_I37 (.Y(N118), .A(N1170), .B(N1171));
NOR2XL inst_cellmath__60_0_I38 (.Y(N120), .A(N1170), .B(N1172));
NOR2XL inst_cellmath__60_0_I39 (.Y(N122), .A(N1170), .B(N1183));
NOR2XL inst_cellmath__60_0_I40 (.Y(N124), .A(N1170), .B(N1184));
NOR2XL inst_cellmath__60_0_I41 (.Y(N126), .A(N1170), .B(N1190));
NOR2XL inst_cellmath__60_0_I42 (.Y(N128), .A(N1170), .B(N1191));
NOR2XL inst_cellmath__60_0_I43 (.Y(N130), .A(N1170), .B(N1192));
NOR2XL inst_cellmath__60_0_I44 (.Y(N132), .A(N1170), .B(N1193));
NOR2XL inst_cellmath__60_0_I45 (.Y(N134), .A(N1170), .B(N1194));
NOR2XL inst_cellmath__60_0_I46 (.Y(N136), .A(N1170), .B(N1195));
OR2XL inst_cellmath__60_0_I47 (.Y(N405), .A(N1170), .B(N1196));
INVXL inst_cellmath__60_0_I52 (.Y(N150), .A(N1171));
NOR2XL inst_cellmath__60_0_I54 (.Y(N154), .A(N1171), .B(N1172));
NOR2XL inst_cellmath__60_0_I55 (.Y(N156), .A(N1171), .B(N1183));
NOR2XL inst_cellmath__60_0_I56 (.Y(N158), .A(N1171), .B(N1184));
NOR2XL inst_cellmath__60_0_I57 (.Y(N160), .A(N1171), .B(N1190));
NOR2XL inst_cellmath__60_0_I58 (.Y(N162), .A(N1171), .B(N1191));
NOR2XL inst_cellmath__60_0_I59 (.Y(N164), .A(N1171), .B(N1192));
NOR2XL inst_cellmath__60_0_I60 (.Y(N166), .A(N1171), .B(N1193));
NOR2XL inst_cellmath__60_0_I61 (.Y(N168), .A(N1171), .B(N1194));
NOR2XL inst_cellmath__60_0_I62 (.Y(N170), .A(N1171), .B(N1195));
OR2XL inst_cellmath__60_0_I63 (.Y(N406), .A(N1171), .B(N1196));
INVXL inst_cellmath__60_0_I68 (.Y(N184), .A(N1172));
NOR2XL inst_cellmath__60_0_I70 (.Y(N188), .A(N1172), .B(N1183));
NOR2XL inst_cellmath__60_0_I71 (.Y(N190), .A(N1172), .B(N1184));
NOR2XL inst_cellmath__60_0_I72 (.Y(N192), .A(N1172), .B(N1190));
NOR2XL inst_cellmath__60_0_I73 (.Y(N194), .A(N1172), .B(N1191));
NOR2XL inst_cellmath__60_0_I74 (.Y(N196), .A(N1172), .B(N1192));
NOR2XL inst_cellmath__60_0_I75 (.Y(N198), .A(N1172), .B(N1193));
NOR2XL inst_cellmath__60_0_I76 (.Y(N200), .A(N1172), .B(N1194));
NOR2XL inst_cellmath__60_0_I77 (.Y(N202), .A(N1172), .B(N1195));
OR2XL inst_cellmath__60_0_I78 (.Y(N407), .A(N1172), .B(N1196));
INVXL inst_cellmath__60_0_I83 (.Y(N216), .A(N1183));
NOR2XL inst_cellmath__60_0_I85 (.Y(N220), .A(N1183), .B(N1184));
NOR2XL inst_cellmath__60_0_I86 (.Y(N222), .A(N1183), .B(N1190));
NOR2XL inst_cellmath__60_0_I87 (.Y(N224), .A(N1183), .B(N1191));
NOR2XL inst_cellmath__60_0_I88 (.Y(N226), .A(N1183), .B(N1192));
NOR2XL inst_cellmath__60_0_I89 (.Y(N228), .A(N1183), .B(N1193));
NOR2XL inst_cellmath__60_0_I90 (.Y(N230), .A(N1183), .B(N1194));
NOR2XL inst_cellmath__60_0_I91 (.Y(N232), .A(N1183), .B(N1195));
OR2XL inst_cellmath__60_0_I92 (.Y(N408), .A(N1183), .B(N1196));
INVXL inst_cellmath__60_0_I97 (.Y(N246), .A(N1184));
NOR2XL inst_cellmath__60_0_I99 (.Y(N250), .A(N1184), .B(N1190));
NOR2XL inst_cellmath__60_0_I100 (.Y(N252), .A(N1184), .B(N1191));
NOR2XL inst_cellmath__60_0_I101 (.Y(N254), .A(N1184), .B(N1192));
NOR2XL inst_cellmath__60_0_I102 (.Y(N256), .A(N1184), .B(N1193));
NOR2XL inst_cellmath__60_0_I103 (.Y(N258), .A(N1184), .B(N1194));
NOR2XL inst_cellmath__60_0_I104 (.Y(N260), .A(N1184), .B(N1195));
OR2XL inst_cellmath__60_0_I105 (.Y(N409), .A(N1184), .B(N1196));
INVXL inst_cellmath__60_0_I110 (.Y(N274), .A(N1190));
NOR2XL inst_cellmath__60_0_I112 (.Y(N278), .A(N1190), .B(N1191));
NOR2XL inst_cellmath__60_0_I113 (.Y(N280), .A(N1190), .B(N1192));
NOR2XL inst_cellmath__60_0_I114 (.Y(N282), .A(N1190), .B(N1193));
NOR2XL inst_cellmath__60_0_I115 (.Y(N284), .A(N1190), .B(N1194));
NOR2XL inst_cellmath__60_0_I116 (.Y(N286), .A(N1190), .B(N1195));
OR2XL inst_cellmath__60_0_I117 (.Y(N410), .A(N1190), .B(N1196));
INVXL inst_cellmath__60_0_I122 (.Y(N300), .A(N1191));
NOR2XL inst_cellmath__60_0_I124 (.Y(N304), .A(N1191), .B(N1192));
NOR2XL inst_cellmath__60_0_I125 (.Y(N306), .A(N1191), .B(N1193));
NOR2XL inst_cellmath__60_0_I126 (.Y(N308), .A(N1191), .B(N1194));
NOR2XL inst_cellmath__60_0_I127 (.Y(N310), .A(N1191), .B(N1195));
OR2XL inst_cellmath__60_0_I128 (.Y(N411), .A(N1191), .B(N1196));
INVXL inst_cellmath__60_0_I133 (.Y(N324), .A(N1192));
NOR2XL inst_cellmath__60_0_I135 (.Y(N328), .A(N1192), .B(N1193));
NOR2XL inst_cellmath__60_0_I136 (.Y(N330), .A(N1192), .B(N1194));
NOR2XL inst_cellmath__60_0_I137 (.Y(N332), .A(N1192), .B(N1195));
OR2XL inst_cellmath__60_0_I138 (.Y(N412), .A(N1192), .B(N1196));
INVXL inst_cellmath__60_0_I143 (.Y(N346), .A(N1193));
NOR2XL inst_cellmath__60_0_I145 (.Y(N350), .A(N1193), .B(N1194));
NOR2XL inst_cellmath__60_0_I146 (.Y(N352), .A(N1193), .B(N1195));
OR2XL inst_cellmath__60_0_I147 (.Y(N413), .A(N1193), .B(N1196));
INVXL inst_cellmath__60_0_I152 (.Y(N366), .A(N1194));
NOR2XL inst_cellmath__60_0_I154 (.Y(N370), .A(N1194), .B(N1195));
OR2XL inst_cellmath__60_0_I155 (.Y(N414), .A(N1194), .B(N1196));
INVXL inst_cellmath__60_0_I160 (.Y(N384), .A(N1195));
ADDHX1 inst_cellmath__60_0_I179 (.CO(N416), .S(N415), .A(N150), .B(N84));
ADDHX1 inst_cellmath__60_0_I180 (.CO(N418), .S(N417), .A(N120), .B(N86));
ADDHX1 inst_cellmath__60_0_I181 (.CO(N420), .S(N419), .A(N184), .B(N88));
ADDFX1 inst_cellmath__60_0_I182 (.CO(N422), .S(N421), .A(N122), .B(N154), .CI(N418));
ADDHX1 inst_cellmath__60_0_I183 (.CO(N424), .S(N423), .A(N156), .B(N90));
ADDFX1 inst_cellmath__60_0_I184 (.CO(N426), .S(N425), .A(N420), .B(N124), .CI(N423));
ADDHX1 inst_cellmath__60_0_I185 (.CO(N428), .S(N427), .A(N216), .B(N92));
ADDFX1 inst_cellmath__60_0_I186 (.CO(N430), .S(N429), .A(N126), .B(N188), .CI(N158));
ADDFX1 inst_cellmath__60_0_I187 (.CO(N432), .S(N431), .A(N427), .B(N424), .CI(N429));
ADDHX1 inst_cellmath__60_0_I188 (.CO(N434), .S(N433), .A(N190), .B(N94));
ADDFX1 inst_cellmath__60_0_I189 (.CO(N436), .S(N435), .A(N128), .B(N160), .CI(N428));
ADDFX1 inst_cellmath__60_0_I190 (.CO(N438), .S(N437), .A(N430), .B(N433), .CI(N435));
ADDHX1 inst_cellmath__60_0_I191 (.CO(N440), .S(N439), .A(N246), .B(N96));
ADDFX1 inst_cellmath__60_0_I192 (.CO(N442), .S(N441), .A(N130), .B(N220), .CI(N162));
ADDFX1 inst_cellmath__60_0_I193 (.CO(N444), .S(N443), .A(N434), .B(N192), .CI(N439));
ADDFX1 inst_cellmath__60_0_I194 (.CO(N446), .S(N445), .A(N441), .B(N436), .CI(N443));
ADDHX1 inst_cellmath__60_0_I195 (.CO(N448), .S(N447), .A(N222), .B(N98));
ADDFX1 inst_cellmath__60_0_I196 (.CO(N450), .S(N449), .A(N132), .B(N194), .CI(N164));
ADDFX1 inst_cellmath__60_0_I197 (.CO(N452), .S(N451), .A(N447), .B(N440), .CI(N442));
ADDFX1 inst_cellmath__60_0_I198 (.CO(N454), .S(N453), .A(N444), .B(N449), .CI(N451));
ADDHX1 inst_cellmath__60_0_I199 (.CO(N456), .S(N455), .A(N274), .B(N100));
ADDFX1 inst_cellmath__60_0_I200 (.CO(N458), .S(N457), .A(N134), .B(N250), .CI(N166));
ADDFX1 inst_cellmath__60_0_I201 (.CO(N460), .S(N459), .A(N196), .B(N224), .CI(N448));
ADDFX1 inst_cellmath__60_0_I202 (.CO(N462), .S(N461), .A(N450), .B(N455), .CI(N457));
ADDFX1 inst_cellmath__60_0_I203 (.CO(N464), .S(N463), .A(N452), .B(N459), .CI(N461));
XNOR2X1 hap1_A_I721 (.Y(N465), .A(N252), .B(N136));
OR2XL hap1_A_I722 (.Y(N466), .A(N252), .B(N136));
ADDFX1 inst_cellmath__60_0_I205 (.CO(N470), .S(N469), .A(N168), .B(N226), .CI(N198));
ADDFX1 inst_cellmath__60_0_I206 (.CO(N472), .S(N471), .A(N456), .B(N404), .CI(N465));
ADDFX1 inst_cellmath__60_0_I207 (.CO(N474), .S(N473), .A(N460), .B(N458), .CI(N469));
ADDFX1 inst_cellmath__60_0_I208 (.CO(N476), .S(N475), .A(N462), .B(N471), .CI(N473));
ADDFX1 inst_cellmath__60_0_I209 (.CO(N478), .S(N477), .A(N278), .B(N300), .CI(N170));
ADDFX1 inst_cellmath__60_0_I210 (.CO(N480), .S(N479), .A(N200), .B(N254), .CI(N228));
ADDFX1 inst_cellmath__60_0_I211 (.CO(N482), .S(N481), .A(N466), .B(N405), .CI(N470));
ADDFX1 inst_cellmath__60_0_I212 (.CO(N484), .S(N483), .A(N479), .B(N477), .CI(N472));
ADDFX1 inst_cellmath__60_0_I213 (.CO(N486), .S(N485), .A(N474), .B(N481), .CI(N483));
ADDFX1 inst_cellmath__60_0_I214 (.CO(N488), .S(N487), .A(N202), .B(N280), .CI(N230));
ADDFX1 inst_cellmath__60_0_I215 (.CO(N490), .S(N489), .A(N406), .B(N256), .CI(N478));
ADDFX1 inst_cellmath__60_0_I216 (.CO(N492), .S(N491), .A(N487), .B(N480), .CI(N482));
ADDFX1 inst_cellmath__60_0_I217 (.CO(N494), .S(N493), .A(N484), .B(N489), .CI(N491));
ADDFX1 inst_cellmath__60_0_I218 (.CO(N496), .S(N495), .A(N304), .B(N324), .CI(N232));
ADDFX1 inst_cellmath__60_0_I219 (.CO(N498), .S(N497), .A(N258), .B(N282), .CI(N407));
ADDFX1 inst_cellmath__60_0_I220 (.CO(N500), .S(N499), .A(N495), .B(N488), .CI(N497));
ADDFX1 inst_cellmath__60_0_I221 (.CO(N502), .S(N501), .A(N492), .B(N490), .CI(N499));
ADDFX1 inst_cellmath__60_0_I222 (.CO(N504), .S(N503), .A(N260), .B(N306), .CI(N284));
ADDFX1 inst_cellmath__60_0_I223 (.CO(N506), .S(N505), .A(N496), .B(N408), .CI(N498));
ADDFX1 inst_cellmath__60_0_I224 (.CO(N508), .S(N507), .A(N500), .B(N503), .CI(N505));
ADDFX1 inst_cellmath__60_0_I225 (.CO(N510), .S(N509), .A(N328), .B(N346), .CI(N286));
ADDFX1 inst_cellmath__60_0_I226 (.CO(N512), .S(N511), .A(N409), .B(N308), .CI(N504));
ADDFX1 inst_cellmath__60_0_I227 (.CO(N514), .S(N513), .A(N506), .B(N509), .CI(N511));
ADDFX1 inst_cellmath__60_0_I228 (.CO(N516), .S(N515), .A(N310), .B(N330), .CI(N410));
ADDFX1 inst_cellmath__60_0_I229 (.CO(N518), .S(N517), .A(N515), .B(N510), .CI(N512));
ADDFX1 inst_cellmath__60_0_I230 (.CO(N520), .S(N519), .A(N350), .B(N366), .CI(N332));
ADDFX1 inst_cellmath__60_0_I231 (.CO(N522), .S(N521), .A(N516), .B(N411), .CI(N519));
ADDFX1 inst_cellmath__60_0_I232 (.CO(N524), .S(N523), .A(N412), .B(N352), .CI(N520));
ADDFX1 inst_cellmath__60_0_I233 (.CO(N526), .S(N525), .A(N370), .B(N384), .CI(N413));
NOR2XL inst_cellmath__60_0_I234 (.Y(N527), .A(N1170), .B(N80));
NOR2XL inst_cellmath__60_0_I236 (.Y(N529), .A(N118), .B(N415));
NAND2XL inst_cellmath__60_0_I237 (.Y(N530), .A(N118), .B(N415));
NOR2XL inst_cellmath__60_0_I238 (.Y(N531), .A(N416), .B(N417));
NAND2XL inst_cellmath__60_0_I239 (.Y(N532), .A(N416), .B(N417));
NOR2XL inst_cellmath__60_0_I240 (.Y(N533), .A(N419), .B(N421));
NAND2XL inst_cellmath__60_0_I241 (.Y(N534), .A(N419), .B(N421));
NOR2XL inst_cellmath__60_0_I242 (.Y(N535), .A(N422), .B(N425));
NAND2XL inst_cellmath__60_0_I243 (.Y(N536), .A(N422), .B(N425));
NOR2XL inst_cellmath__60_0_I244 (.Y(N537), .A(N426), .B(N431));
NAND2XL inst_cellmath__60_0_I245 (.Y(N538), .A(N426), .B(N431));
AND2XL inst_cellmath__60_0_I248 (.Y(N541), .A(N528), .B(N527));
INVXL inst_cellmath__60_0_I794 (.Y(N1203), .A(N529));
INVXL inst_cellmath__60_0_I795 (.Y(N1204), .A(N530));
OAI21XL inst_cellmath__60_0_I256 (.Y(N551), .A0(N1204), .A1(N541), .B0(N1203));
AOI21XL inst_cellmath__60_0_I264 (.Y(N559), .A0(N532), .A1(N551), .B0(N531));
INVXL inst_cellmath__60_0_I801 (.Y(N1210), .A(N533));
INVXL inst_cellmath__60_0_I802 (.Y(N1211), .A(N534));
OAI21XL inst_cellmath__60_0_I276 (.Y(N571), .A0(N1211), .A1(N559), .B0(N1210));
AOI21XL inst_cellmath__60_0_I288 (.Y(N583), .A0(N536), .A1(N571), .B0(N535));
INVXL inst_cellmath__60_0_I812 (.Y(N1221), .A(N537));
INVXL inst_cellmath__60_0_I813 (.Y(N1222), .A(N538));
OAI21XL inst_cellmath__60_0_I304 (.Y(N632), .A0(N1222), .A1(N583), .B0(N1221));
NAND2BXL inst_cellmath__60_0_I314 (.Y(N611), .AN(N529), .B(N530));
NAND2BXL inst_cellmath__60_0_I317 (.Y(N614), .AN(N531), .B(N532));
NAND2BXL inst_cellmath__60_0_I320 (.Y(N617), .AN(N533), .B(N534));
NAND2BXL inst_cellmath__60_0_I323 (.Y(N620), .AN(N535), .B(N536));
NAND2BXL inst_cellmath__60_0_I326 (.Y(N623), .AN(N537), .B(N538));
XOR2XL inst_cellmath__60_0_I1367 (.Y(inst_cellmath__60_0_out0[2]), .A(N1170), .B(N80));
XOR2XL inst_cellmath__60_0_I828 (.Y(inst_cellmath__60_0_out0[3]), .A(N527), .B(N528));
XNOR2X1 inst_cellmath__60_0_I822 (.Y(inst_cellmath__60_0_out0[4]), .A(N541), .B(N611));
XOR2XL inst_cellmath__60_0_I829 (.Y(inst_cellmath__60_0_out0[5]), .A(N551), .B(N614));
XNOR2X1 inst_cellmath__60_0_I836 (.Y(inst_cellmath__60_0_out0[6]), .A(N559), .B(N617));
XOR2XL inst_cellmath__60_0_I825 (.Y(inst_cellmath__60_0_out0[7]), .A(N571), .B(N620));
XNOR2X1 inst_cellmath__60_0_I333 (.Y(inst_cellmath__60_0_out0[8]), .A(N583), .B(N623));
NOR2XL inst_cellmath__60_0_I336 (.Y(N634), .A(N432), .B(N437));
XOR2XL inst_cellmath__60_0_I337 (.Y(N635), .A(N432), .B(N437));
NOR2XL inst_cellmath__60_0_I338 (.Y(N636), .A(N438), .B(N445));
XOR2XL inst_cellmath__60_0_I339 (.Y(N637), .A(N438), .B(N445));
NOR2XL inst_cellmath__60_0_I340 (.Y(N638), .A(N446), .B(N453));
XOR2XL inst_cellmath__60_0_I341 (.Y(N639), .A(N446), .B(N453));
NOR2XL inst_cellmath__60_0_I342 (.Y(N640), .A(N454), .B(N463));
XOR2XL inst_cellmath__60_0_I343 (.Y(N641), .A(N454), .B(N463));
NOR2XL inst_cellmath__60_0_I344 (.Y(N642), .A(N464), .B(N475));
XOR2XL inst_cellmath__60_0_I345 (.Y(N643), .A(N464), .B(N475));
NOR2XL inst_cellmath__60_0_I346 (.Y(N644), .A(N476), .B(N485));
XOR2XL inst_cellmath__60_0_I347 (.Y(N645), .A(N476), .B(N485));
NOR2XL inst_cellmath__60_0_I348 (.Y(N646), .A(N486), .B(N493));
XOR2XL inst_cellmath__60_0_I349 (.Y(N647), .A(N486), .B(N493));
NOR2XL inst_cellmath__60_0_I350 (.Y(N648), .A(N494), .B(N501));
XOR2XL inst_cellmath__60_0_I351 (.Y(N649), .A(N494), .B(N501));
NOR2XL inst_cellmath__60_0_I352 (.Y(N650), .A(N502), .B(N507));
XOR2XL inst_cellmath__60_0_I353 (.Y(N651), .A(N502), .B(N507));
NOR2XL inst_cellmath__60_0_I354 (.Y(N652), .A(N508), .B(N513));
XOR2XL inst_cellmath__60_0_I355 (.Y(N653), .A(N508), .B(N513));
NOR2XL inst_cellmath__60_0_I356 (.Y(N654), .A(N517), .B(N514));
XOR2XL inst_cellmath__60_0_I357 (.Y(N655), .A(N517), .B(N514));
NOR2XL inst_cellmath__60_0_I358 (.Y(N656), .A(N518), .B(N521));
XOR2XL inst_cellmath__60_0_I359 (.Y(N657), .A(N518), .B(N521));
NOR2XL inst_cellmath__60_0_I360 (.Y(N658), .A(N523), .B(N522));
XOR2XL inst_cellmath__60_0_I361 (.Y(N659), .A(N523), .B(N522));
NOR2XL inst_cellmath__60_0_I362 (.Y(N660), .A(N525), .B(N524));
XOR2XL inst_cellmath__60_0_I363 (.Y(N661), .A(N525), .B(N524));
NOR2XL inst_cellmath__60_0_I364 (.Y(N662), .A(N414), .B(N526));
XOR2XL inst_cellmath__60_0_I365 (.Y(N663), .A(N414), .B(N526));
NAND2BXL inst_cellmath__60_0_I748 (.Y(N665), .AN(N1196), .B(N1195));
AO21XL inst_cellmath__60_0_I370 (.Y(N668), .A0(N635), .A1(N632), .B0(N634));
AO21XL inst_cellmath__60_0_I376 (.Y(N674), .A0(N637), .A1(N668), .B0(N636));
AO21XL inst_cellmath__60_0_I384 (.Y(N682), .A0(N639), .A1(N674), .B0(N638));
AO21XL inst_cellmath__60_0_I394 (.Y(N692), .A0(N641), .A1(N682), .B0(N640));
AO21XL inst_cellmath__60_0_I406 (.Y(N704), .A0(N643), .A1(N692), .B0(N642));
AO21XL inst_cellmath__60_0_I420 (.Y(N718), .A0(N645), .A1(N704), .B0(N644));
AO21XL inst_cellmath__60_0_I436 (.Y(N734), .A0(N647), .A1(N718), .B0(N646));
AO21XL inst_cellmath__60_0_I454 (.Y(N752), .A0(N649), .A1(N734), .B0(N648));
AO21XL inst_cellmath__60_0_I474 (.Y(N772), .A0(N651), .A1(N752), .B0(N650));
AO21XL inst_cellmath__60_0_I496 (.Y(N794), .A0(N653), .A1(N772), .B0(N652));
AO21XL inst_cellmath__60_0_I520 (.Y(N818), .A0(N655), .A1(N794), .B0(N654));
AO21XL inst_cellmath__60_0_I546 (.Y(N844), .A0(N657), .A1(N818), .B0(N656));
AO21XL inst_cellmath__60_0_I574 (.Y(N872), .A0(N659), .A1(N844), .B0(N658));
AO21XL inst_cellmath__60_0_I604 (.Y(N902), .A0(N661), .A1(N872), .B0(N660));
AO21XL inst_cellmath__60_0_I636 (.Y(N934), .A0(N663), .A1(N902), .B0(N662));
XNOR2X1 inst_cellmath__60_0_I676 (.Y(inst_cellmath__60_0_out0[9]), .A(N632), .B(N635));
XNOR2X1 inst_cellmath__60_0_I749 (.Y(inst_cellmath__60_0_out0[10]), .A(N668), .B(N637));
XNOR2X1 inst_cellmath__60_0_I1368 (.Y(inst_cellmath__60_0_out0[11]), .A(N674), .B(N639));
XNOR2X1 inst_cellmath__60_0_I679 (.Y(inst_cellmath__60_0_out0[12]), .A(N682), .B(N641));
XNOR2X1 inst_cellmath__60_0_I680 (.Y(inst_cellmath__60_0_out0[13]), .A(N692), .B(N643));
XNOR2X1 inst_cellmath__60_0_I681 (.Y(inst_cellmath__60_0_out0[14]), .A(N704), .B(N645));
XNOR2X1 inst_cellmath__60_0_I682 (.Y(inst_cellmath__60_0_out0[15]), .A(N718), .B(N647));
XNOR2X1 inst_cellmath__60_0_I683 (.Y(inst_cellmath__60_0_out0[16]), .A(N734), .B(N649));
XNOR2X1 inst_cellmath__60_0_I684 (.Y(inst_cellmath__60_0_out0[17]), .A(N752), .B(N651));
XNOR2X1 inst_cellmath__60_0_I685 (.Y(inst_cellmath__60_0_out0[18]), .A(N772), .B(N653));
XNOR2X1 inst_cellmath__60_0_I686 (.Y(inst_cellmath__60_0_out0[19]), .A(N794), .B(N655));
XNOR2X1 inst_cellmath__60_0_I687 (.Y(inst_cellmath__60_0_out0[20]), .A(N818), .B(N657));
XNOR2X1 inst_cellmath__60_0_I688 (.Y(inst_cellmath__60_0_out0[21]), .A(N844), .B(N659));
XNOR2X1 inst_cellmath__60_0_I689 (.Y(inst_cellmath__60_0_out0[22]), .A(N872), .B(N661));
XNOR2X1 inst_cellmath__60_0_I690 (.Y(inst_cellmath__60_0_out0[23]), .A(N902), .B(N663));
XNOR2X1 inst_cellmath__60_0_I691 (.Y(inst_cellmath__60_0_out0[24]), .A(N934), .B(N665));
assign inst_cellmath__60_0_out0[0] = inst_cellmath__60_0_in1[3];
assign inst_cellmath__60_0_out0[1] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_noninc_a_cellmath__55_2WWMM_bdw1412651405_bdw (
	inst_noninc_a_cellmath__55_2WWMM_out0,
	inst_noninc_a_cellmath__55_2WWMM_in0
	); /* architecture "gate_level" */ 
output [52:0] inst_noninc_a_cellmath__55_2WWMM_out0;
input [22:16] inst_noninc_a_cellmath__55_2WWMM_in0;
wire N1044,N1045,N1060,N1061,N1062,N1066,N1068 
	,N1084,N1086,N1089,N1092,N1093,N1102,N1103,N2138 
	,N2140,N2141,N2142,N2146,N2147,N2163,N2166,N2168 
	,N2170,N2174,N2175,N2176,N2179,N2180,N2199,N2200 
	,N2201,N2202,N2203,N2211,N2212,N2213,N2214,N2215 
	,N2216,N2217,N2218,N2219,N2220,N2221,N2222,N2223 
	,N2236,N2237,N2238,N2239,N2240,N2241,N2242,N2243 
	,N2244,N2245,N2246,N2247,N2248,N2249,N2250,N2251 
	,N2253,N2256,N2257,N2258,N2259,N2261,N3281,N3282 
	,N3287,N3304,N3305,N3306,N3309,N3314,N3322,N3327 
	,N4329,N4342,N4344,N4345,N4346,N4350,N4351,N4367 
	,N4371,N4376,N4377,N4380,N4382,N4396,N4411,N4413 
	,N4414,N4415,N4416,N4417,N4425,N4426,N4427,N4428 
	,N4429,N4430,N4431,N4432,N4433,N4434,N4435,N4436 
	,N4437,N4448,N4449,N4450,N4451,N4452,N4453,N4454 
	,N4455,N4456,N4457,N4458,N4459,N4461,N4462,N4463 
	,N4464,N4465,N4466,N4467,N4468,N4469,N4470,N4473 
	,N4478,N4479,N4480,N4481,N4482,N4483,N4493,N4494 
	,N4495,N4496,N4497,N4498,N4499,N4500,N4501,N4502 
	,N4503,N4504,N4505,N4506,N4507,N4513,N4514,N4515 
	,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4523 
	,N4524,N4525,N4526,N4527,N4528,N4529,N4530,N4531 
	,N4532,N4533,N4534,N4535,N5537,N5550,N5553,N5554 
	,N5555,N5558,N5578,N5584,N5586,N5591,N5592,N5593 
	,N5594,N6610,N6613,N6633,N6635,N6638,N6641,N6642 
	,N6643,N6648,N6657,N6670,N6671,N6672,N6673,N6683 
	,N6684,N6685,N6686,N6687,N6690,N6691,N6692,N6693 
	,N6694,N6695,N6696,N6697,N6698,N6707,N6708,N6709 
	,N6710,N6711,N6712,N6713,N6714,N6715,N6716,N6717 
	,N6718,N6719,N6720,N6721,N6722,N6723,N6724,N6725 
	,N6726,N6727,N7736,N7739,N7753,N7755,N7759,N7780 
	,N7783,N7790,N7795,N7799,N8814,N8819,N8831,N8843 
	,N8845,N8861,N8862,N8863,N8867,N8868,N8870,N8871 
	,N8873,N8895,N8896,N8897,N8898,N8899,N8900,N8901 
	,N8909,N8910,N8911,N8912,N8913,N8914,N8915,N8916 
	,N8917,N8919,N8922,N8923,N8924,N8925,N8926,N8933 
	,N8934,N8935,N8936,N8937,N8938,N8939,N8940,N8941 
	,N8942,N8943,N8944,N8945,N8946,N8947,N8948,N8949 
	,N8950,N8951,N8952,N8953,N8954,N8962,N8963,N8964 
	,N8965,N8966,N8967,N8968,N8972,N8977,N8978,N8979 
	,N8980,N8981,N8982,N8983,N8984,N8985,N8986,N8987 
	,N8988,N8989,N8990,N8991,N8998,N8999,N9000,N9001 
	,N9002,N9003,N9004,N9005,N9006,N9007,N9008,N9009 
	,N9010,N9011,N9012,N9013,N9014,N9015,N9016,N9017 
	,N9018,N9019,N9020,N9022,N9028,N9029,N9030,N9031 
	,N9032,N9033,N9034,N9036,N9039,N9042,N9043,N9044 
	,N9045,N9046,N9047,N9048,N9049,N9050,N9051,N9052 
	,N9053,N9054,N9055,N9056,N9057,N9063,N9064,N9065 
	,N9066,N9067,N9068,N9069,N9070,N9071,N9072,N9073 
	,N9074,N9075,N9076,N9077,N9078,N9079,N9080,N9081 
	,N9082,N9083,N9084,N9085,N9086,N10112,N10134,N10137 
	,N10146,N11159,N11176,N11178,N11181,N11204,N11207,N11210 
	,N11236,N11237,N11238,N11239,N11240,N11241,N11242,N11243 
	,N11248,N11249,N11250,N11251,N11252,N11253,N11254,N11255 
	,N11256,N11257,N11258,N11259,N11271,N11272,N11273,N11274 
	,N11275,N11276,N11277,N11278,N11279,N11280,N11281,N11282 
	,N11283,N11284,N11285,N11286,N11287,N11292,N11293,N11294 
	,N11295,N11296,N12316,N12319,N12328,N12343,N12346,N12357 
	,N12362,N12363,N12366,N12367,N13404,N13406,N13407,N13408 
	,N13411,N13437,N13443,N13448,N13459,N13462,N13471,N13472 
	,N13473,N13476,N13477,N13478,N13487,N13488,N13489,N13490 
	,N13491,N13492,N13493,N13494,N13495,N13496,N13497,N13498 
	,N13499,N13501,N13508,N13509,N13510,N13511,N13512,N13513 
	,N13514,N13515,N13516,N13517,N13518,N13519,N13520,N13521 
	,N13522,N13523,N13524,N13525,N13526,N13527,N13528,N13529 
	,N13538,N13539,N13540,N13541,N13542,N13543,N13544,N13545 
	,N13546,N13551,N13552,N13553,N13554,N13555,N13556,N13557 
	,N13558,N13559,N13560,N13561,N13562,N13563,N13564,N13565 
	,N13566,N13567,N13569,N13572,N13573,N13574,N13575,N13576 
	,N13577,N13578,N13579,N13580,N13581,N13582,N13583,N13584 
	,N13585,N13586,N13587,N13588,N13589,N13590,N13591,N13592 
	,N13593,N13594,N14617,N14619,N14621,N14638,N14641,N14649 
	,N14658,N15695,N15708,N15724,N15725,N15750,N15751,N15752 
	,N15753,N15754,N15755,N15756,N15762,N15763,N15764,N15765 
	,N15766,N15767,N15768,N15769,N15770,N15771,N15772,N15773 
	,N15774,N15775,N15776,N15783,N15784,N15785,N15786,N15787 
	,N15788,N15789,N15790,N15791,N15792,N15793,N15794,N15795 
	,N15796,N15797,N15798,N15799,N15800,N15801,N15802,N15804 
	,N15805,N16832,N16845,N16861,N16862,N16869,N16878,N16879 
	,N16882,N17901,N17908,N17948,N17951,N17969,N17970,N17971 
	,N17972,N17973,N17974,N17975,N17976,N17982,N17983,N17984 
	,N17985,N17986,N17987,N17989,N17990,N17991,N17992,N17993 
	,N17994,N17995,N17996,N17997,N17998,N18002,N18003,N18004 
	,N18005,N18006,N18007,N18008,N18009,N18010,N18011,N18012 
	,N18013,N18014,N18015,N18016,N18017,N18018,N18019,N18020 
	,N18023,N18024,N18025,N18026,N18034,N18035,N18036,N18037 
	,N18038,N18039,N18040,N18041,N18046,N18047,N18048,N18049 
	,N18050,N18051,N18052,N18053,N18054,N18055,N18056,N18057 
	,N18058,N18059,N18060,N18061,N18062,N18067,N18068,N18069 
	,N18070,N18071,N18072,N18073,N18074,N18075,N18076,N18077 
	,N18078,N18079,N18080,N18081,N18082,N18083,N18084,N18085 
	,N18086,N18087,N18088,N18089,N18090,N18094,N18095,N18096 
	,N18097,N18098,N18099,N18100,N18101,N18102,N18103,N18106 
	,N18107,N18108,N18109,N18110,N18111,N18112,N18113,N18114 
	,N18115,N18116,N18117,N18118,N18119,N18120,N18121,N18122 
	,N18125,N18126,N18127,N18128,N18129,N18130,N18131,N18132 
	,N18133,N18134,N18135,N18136,N18137,N18138,N18139,N18140 
	,N18141,N18142,N18143,N18144,N18145,N18146,N18147,N18148 
	,N18215,N18217,N18219,N18221,N18223,N18225,N18227,N18229 
	,N18231,N18233,N18235,N18239,N18241,N18243,N18245,N18247 
	,N18253,N18255,N18257,N18259,N18261,N18265,N18267,N18269 
	,N18271,N18273,N18275,N18277,N18279,N18281,N18283,N18285 
	,N18287,N18289,N18291,N18293,N18295,N18297,N18299,N18301 
	,N18303,N18305,N18307,N18309,N18311,N18313,N18315,N18317 
	,N18319,N18321,N18323,N18325,N18327,N18329,N18331,N18333 
	,N18335,N18337,N18339,N18341,N18343,N18345,N18347,N18349 
	,N18351,N18353,N18355,N18357,N18359,N18361,N18405,N18416 
	,N18424,N18544,N18557,N18581,N18589,N18607,N18714,N18818 
	,N18881,N18896,N18972,N19053,N19055,N19150,N19157,N19164 
	,N19171,N19178;
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13734 (.Y(N18405), .A(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I13745 (.Y(N18416), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I14498 (.Y(N18424), .A0(N18405), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I323 (.Y(N18215), .A(N18416), .B(N18405));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I333 (.Y(N18217), .A(N18416), .B(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I334 (.Y(N18219), .A(N18416), .B(N18405));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I339 (.Y(N18221), .A(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I696 (.Y(N18223), .A(N18416), .B(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I727 (.Y(N18225), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I731 (.Y(N18227), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B(N18405));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I13873 (.Y(N18544), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I749 (.Y(N18229), .A0(N18544), .A1(N18215), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I750 (.Y(N1044), .A0(N18544), .A1(N18223), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I751 (.Y(N1045), .A0(N18544), .A1(N18221), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I752 (.Y(N18231), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18219));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I759 (.Y(N1060), .A0(N18544), .A1(N18219), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I760 (.Y(N1061), .A0(N18544), .A1(N18416), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I761 (.Y(N1062), .A(N18217));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I762 (.Y(N18233), .A0(N18544), .A1(N18217), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I763 (.Y(N18235), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13886 (.Y(N18557), .A(N18424));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I765 (.Y(N1066), .A0(N18544), .A1(N18223), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I766 (.Y(N18239), .A0(N18544), .A1(N18416), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I767 (.Y(N1068), .A(N18544), .B(N18221));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I777 (.Y(N1084), .A0(N18544), .A1(N18223), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I779 (.Y(N1086), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I780 (.Y(N18241), .A0(N18544), .A1(N18221), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I781 (.Y(N18243), .A0(N18544), .A1(N18225), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I782 (.Y(N1089), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18223));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I783 (.Y(N1092), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I784 (.Y(N1093), .A(N18544), .B(N18219));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I785 (.Y(N18245), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18227));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I786 (.Y(N18247), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I788 (.Y(N1102), .A0(N18544), .A1(N18416), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I789 (.Y(N1103), .A0(N18544), .A1(N18219), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I14481 (.Y(N18581), .A(N18405), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I14499 (.Y(N18589), .A0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18416), .B1(N18405));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1551 (.Y(N18253), .A(N18544), .B(N18225));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1554 (.Y(N18255), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1555 (.Y(N18257), .A(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1561 (.Y(N18259), .A0(N18544), .A1(N18589), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1562 (.Y(N2138), .A(N18544), .B(N18405));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1563 (.Y(N2140), .A0(N18544), .A1(N18424), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1564 (.Y(N2141), .A0(N18544), .A1(N18221), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1565 (.Y(N2142), .A0(N18544), .A1(N18219), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1566 (.Y(N18261), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1569 (.Y(N2146), .A0(N18544), .A1(N18589), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1570 (.Y(N2147), .A0(N18544), .A1(N18581), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13936 (.Y(N18607), .A(N18589));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1572 (.Y(N18265), .A0(N18544), .A1(N18215), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1573 (.Y(N18267), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18215));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1574 (.Y(N18269), .A(N18544), .B(N18225));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1580 (.Y(N2163), .A(N18405), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1581 (.Y(N18271), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1582 (.Y(N2166), .A0(N18544), .A1(N18225), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1583 (.Y(N18273), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1584 (.Y(N2168), .A(N18544), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1585 (.Y(N2170), .A(N18544), .B(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1588 (.Y(N2174), .A0(N18544), .A1(N18215), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1589 (.Y(N2175), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1590 (.Y(N2176), .A0(N18544), .A1(N18223), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1592 (.Y(N18275), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1593 (.Y(N2179), .A0(N18544), .A1(N18589), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1594 (.Y(N2180), .A0(N18544), .A1(N18219), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1596 (.Y(N18277), .A0(N18544), .A1(N18405), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1597 (.Y(N18279), .A0(N18544), .A1(N18424), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1598 (.Y(N18281), .A0(N18544), .A1(N18225), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I14301 (.Y(N18972), .A(inst_noninc_a_cellmath__55_2WWMM_in0[19]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14384 (.Y(N19055), .A(N18972));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I14043 (.Y(N18714), .A(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1605 (.Y(N2199), .A0(N18714), .A1(N18253), .B0(N18229), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1606 (.Y(N2200), .A0(N18714), .A1(N18405), .B0(N1044), .B1(N19055));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14382 (.Y(N19053), .A(N18972));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1607 (.Y(N2201), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N1045), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1608 (.Y(N2202), .A0(N18714), .A1(N18255), .B0(N18231), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1609 (.Y(N2203), .A(N18714), .B(N18257));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1615 (.Y(N2211), .A0(N18714), .A1(N18259), .B0(N1060), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1616 (.Y(N2212), .A0(N18714), .A1(N2138), .B0(N1061), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1617 (.Y(N2213), .A0(N18714), .A1(N2140), .B0(N1062), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1618 (.Y(N2214), .A0(N18714), .A1(N2141), .B0(N18233), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1619 (.Y(N2215), .A0(N18714), .A1(N2142), .B0(N18235), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1620 (.Y(N2216), .A0(N18714), .A1(N18261), .B0(N18557), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1621 (.Y(N2217), .A0(N18714), .A1(N18235), .B0(N1066), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1622 (.Y(N2218), .A0(N18714), .A1(N18261), .B0(N18239), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1623 (.Y(N2219), .A0(N18714), .A1(N2146), .B0(N1068), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1624 (.Y(N2220), .A0(N18714), .A1(N2147), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1625 (.Y(N2221), .A0(N18714), .A1(N18607), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1626 (.Y(N2222), .A0(N18714), .A1(N18265), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1627 (.Y(N2223), .A(N19055), .B(N18267));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1628 (.Y(N18283), .A(N19053), .B(N18269));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1633 (.Y(N2236), .A0(N18714), .A1(N18247), .B0(N1084), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1634 (.Y(N2237), .A0(N18714), .A1(N2163), .B0(N18233), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1635 (.Y(N2238), .A0(N18714), .A1(N18271), .B0(N1086), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1636 (.Y(N2239), .A0(N18714), .A1(N2166), .B0(N18241), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1637 (.Y(N2240), .A0(N18714), .A1(N18273), .B0(N18243), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1638 (.Y(N2241), .A0(N18714), .A1(N2168), .B0(N1089), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1639 (.Y(N2242), .A0(N18714), .A1(N2170), .B0(N1092), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1640 (.Y(N2243), .A0(N18714), .A1(N18243), .B0(N1093), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1641 (.Y(N2244), .A0(N18714), .A1(N18271), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1642 (.Y(N2245), .A0(N18714), .A1(N2174), .B0(N18247), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1643 (.Y(N2246), .A0(N18714), .A1(N2175), .B0(N18557), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1644 (.Y(N2247), .A0(N18714), .A1(N2176), .B0(N1102), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1645 (.Y(N2248), .A0(N18714), .A1(N18273), .B0(N1103), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1646 (.Y(N2249), .A0(N18714), .A1(N18275), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1647 (.Y(N2250), .A0(N18714), .A1(N2179), .B0(N18247), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1648 (.Y(N2251), .A(N18714), .B(N2180));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1649 (.Y(N2253), .A(N19053), .B(N18253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1650 (.Y(N2256), .A0(N18714), .A1(N18277), .B0(N18405), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1651 (.Y(N2257), .A0(N18714), .A1(N18279), .B0(N18416), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1652 (.Y(N2258), .A0(N18714), .A1(N18281), .B0(N18544), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1653 (.Y(N2259), .A(N18714), .B(N18269));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1654 (.Y(N2261), .A(N18714), .B(N18267));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2411 (.Y(N18285), .A(N18544), .B(N18416));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2417 (.Y(N18287), .A0(N18544), .A1(N18215), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2418 (.Y(N18289), .A0(N18544), .A1(N18223), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2419 (.Y(N3281), .A0(N18544), .A1(N18221), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2420 (.Y(N3282), .A0(N18544), .A1(N18225), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2423 (.Y(N3287), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18225));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2424 (.Y(N18291), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2425 (.Y(N18293), .A0(N18544), .A1(N18589), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2426 (.Y(N18295), .A0(N18544), .A1(N18581), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2427 (.Y(N18297), .A0(N18544), .A1(N18424), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2428 (.Y(N18299), .A0(N18544), .A1(N18219), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I2429 (.Y(N18301), .A(N18544), .B(N18221));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2435 (.Y(N3304), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2436 (.Y(N3305), .A0(N18544), .A1(N18227), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2437 (.Y(N3306), .A(N18544), .B(N18215));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I2438 (.Y(N3309), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18221));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2440 (.Y(N18303), .A0(N18544), .A1(N18589), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2441 (.Y(N3314), .A0(N18544), .A1(N18581), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2444 (.Y(N18305), .A0(N18544), .A1(N18217), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2448 (.Y(N3322), .A0(N18544), .A1(N18581), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2449 (.Y(N18307), .A0(N18544), .A1(N18219), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2450 (.Y(N18309), .A0(N18544), .A1(N18227), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2452 (.Y(N18311), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2453 (.Y(N3327), .A0(N18544), .A1(N18416), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I2454 (.Y(N18313), .A0(N18544), .A1(N18416), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3210 (.Y(N4329), .A0(N18544), .A1(N18405), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3219 (.Y(N4342), .A0(N18544), .A1(N18219), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3220 (.Y(N18315), .A0(N18544), .A1(N18215), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I3221 (.Y(N4344), .A(N18215));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3222 (.Y(N4345), .A0(N18544), .A1(N18227), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3223 (.Y(N4346), .A(N18225), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3224 (.Y(N18317), .A(N18544), .B(N18581));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3225 (.Y(N4350), .A0(N18544), .A1(N18416), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3226 (.Y(N4351), .A0(N18544), .A1(N18416), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3228 (.Y(N18319), .A0(N18544), .A1(N18223), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3229 (.Y(N18321), .A0(N18544), .A1(N18217), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3231 (.Y(N18323), .A(N18215), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3237 (.Y(N4367), .A(N18544), .B(inst_noninc_a_cellmath__55_2WWMM_in0[16]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3239 (.Y(N4371), .A(N18544), .B(N18217));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3241 (.Y(N4376), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3242 (.Y(N4377), .A0(N18544), .A1(N18219), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3245 (.Y(N4380), .A0(N18544), .A1(N18581), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3247 (.Y(N4382), .A(N18544), .B(N18227));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3248 (.Y(N18325), .A0(N18544), .A1(N18581), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3255 (.Y(N4396), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3256 (.Y(N18327), .A(N18544), .B(N18219));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3263 (.Y(N4411), .A(N18714), .B(N2168));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3264 (.Y(N4413), .A0(N18714), .A1(N4329), .B0(N18405), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3265 (.Y(N4414), .A0(N18714), .A1(N18293), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3266 (.Y(N4415), .A0(N18714), .A1(N18299), .B0(N18255), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3267 (.Y(N4416), .A0(N18714), .A1(N18257), .B0(N18285), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3268 (.Y(N4417), .A(N18714), .B(N18257));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3273 (.Y(N4425), .A0(N18714), .A1(N4342), .B0(N18287), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3274 (.Y(N4426), .A0(N18714), .A1(N18315), .B0(N18289), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3275 (.Y(N4427), .A0(N18714), .A1(N4344), .B0(N3281), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3276 (.Y(N4428), .A0(N18714), .A1(N4345), .B0(N3282), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3277 (.Y(N4429), .A0(N18714), .A1(N4346), .B0(N18241), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3278 (.Y(N4430), .A0(N18714), .A1(N18317), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3279 (.Y(N4431), .A0(N18714), .A1(N4350), .B0(N3287), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3280 (.Y(N4432), .A0(N18714), .A1(N4351), .B0(N18291), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3281 (.Y(N4433), .A0(N18714), .A1(N2179), .B0(N18293), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3282 (.Y(N4434), .A0(N18714), .A1(N18319), .B0(N18295), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3283 (.Y(N4435), .A0(N18714), .A1(N18321), .B0(N18297), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3284 (.Y(N4436), .A0(N18714), .A1(N18313), .B0(N18299), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3285 (.Y(N4437), .A0(N18714), .A1(N18323), .B0(N18301), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3286 (.Y(N18329), .A(N18714), .B(N18323));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3291 (.Y(N4448), .A0(N18714), .A1(N4367), .B0(N3304), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3292 (.Y(N4449), .A0(N18714), .A1(N18303), .B0(N3305), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3293 (.Y(N4450), .A0(N18714), .A1(N4371), .B0(N3306), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3294 (.Y(N4451), .A0(N18714), .A1(N18253), .B0(N3309), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3295 (.Y(N4452), .A0(N18714), .A1(N4376), .B0(N18233), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3296 (.Y(N4453), .A0(N18714), .A1(N4377), .B0(N18303), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3297 (.Y(N4454), .A0(N18714), .A1(N2174), .B0(N3314), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3298 (.Y(N4455), .A0(N18714), .A1(N18287), .B0(N18241), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3299 (.Y(N4456), .A0(N18714), .A1(N4380), .B0(N18239), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3300 (.Y(N4457), .A0(N18714), .A1(N18311), .B0(N18305), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3301 (.Y(N4458), .A0(N18714), .A1(N4382), .B0(N18305), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3302 (.Y(N4459), .A(N18714), .B(N18325));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3303 (.Y(N4461), .A0(N18714), .A1(N18229), .B0(N3282), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3304 (.Y(N4462), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N3322), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3305 (.Y(N4463), .A0(N18714), .A1(N18247), .B0(N18307), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3306 (.Y(N4464), .A0(N18714), .A1(N18405), .B0(N18309), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3307 (.Y(N4465), .A0(N18714), .A1(N18416), .B0(N18271), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3308 (.Y(N4466), .A0(N18714), .A1(N18291), .B0(N18311), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3309 (.Y(N4467), .A0(N18714), .A1(N4396), .B0(N3327), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3310 (.Y(N4468), .A0(N18714), .A1(N18327), .B0(N18313), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3311 (.Y(N4469), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B0(N18247), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3312 (.Y(N4470), .A(N19055), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3313 (.Y(N4473), .A(N18714), .B(N18544));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I14147 (.Y(N18818), .A(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3317 (.Y(N4478), .A0(N18818), .A1(N4411), .B0(N2199), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3318 (.Y(N4479), .A0(N18818), .A1(N4413), .B0(N2200), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3319 (.Y(N4480), .A0(N18818), .A1(N4414), .B0(N2201), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3320 (.Y(N4481), .A0(N18818), .A1(N4415), .B0(N2202), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3321 (.Y(N4482), .A0(N18818), .A1(N4416), .B0(N2203), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3322 (.Y(N4483), .A(inst_noninc_a_cellmath__55_2WWMM_in0[20]), .B(N4417));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3327 (.Y(N4493), .A0(N18818), .A1(N4425), .B0(N2211), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3328 (.Y(N4494), .A0(N18818), .A1(N4426), .B0(N2212), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3329 (.Y(N4495), .A0(N18818), .A1(N4427), .B0(N2213), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3330 (.Y(N4496), .A0(N18818), .A1(N4428), .B0(N2214), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3331 (.Y(N4497), .A0(N18818), .A1(N4429), .B0(N2215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3332 (.Y(N4498), .A0(N18818), .A1(N4430), .B0(N2216), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3333 (.Y(N4499), .A0(N18818), .A1(N4431), .B0(N2217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3334 (.Y(N4500), .A0(N18818), .A1(N4432), .B0(N2218), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3335 (.Y(N4501), .A0(N18818), .A1(N4433), .B0(N2219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3336 (.Y(N4502), .A0(N18818), .A1(N4434), .B0(N2220), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3337 (.Y(N4503), .A0(N18818), .A1(N4435), .B0(N2221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3338 (.Y(N4504), .A0(N18818), .A1(N4436), .B0(N2222), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3339 (.Y(N4505), .A0(N18818), .A1(N4437), .B0(N2223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3340 (.Y(N4506), .A0(N18818), .A1(N18329), .B0(N18283), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I3341 (.Y(N4507), .A(N18818), .B(N2253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3345 (.Y(N4513), .A0(N18818), .A1(N4448), .B0(N2236), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3346 (.Y(N4514), .A0(N18818), .A1(N4449), .B0(N2237), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3347 (.Y(N4515), .A0(N18818), .A1(N4450), .B0(N2238), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3348 (.Y(N4516), .A0(N18818), .A1(N4451), .B0(N2239), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3349 (.Y(N4517), .A0(N18818), .A1(N4452), .B0(N2240), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3350 (.Y(N4518), .A0(N18818), .A1(N4453), .B0(N2241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3351 (.Y(N4519), .A0(N18818), .A1(N4454), .B0(N2242), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3352 (.Y(N4520), .A0(N18818), .A1(N4455), .B0(N2243), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3353 (.Y(N4521), .A0(N18818), .A1(N4456), .B0(N2244), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3354 (.Y(N4522), .A0(N18818), .A1(N4457), .B0(N2245), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3355 (.Y(N4523), .A0(N18818), .A1(N4458), .B0(N2246), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3356 (.Y(N4524), .A0(N18818), .A1(N4459), .B0(N2247), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3357 (.Y(N4525), .A0(N18818), .A1(N4461), .B0(N2248), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3358 (.Y(N4526), .A0(N18818), .A1(N4462), .B0(N2249), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3359 (.Y(N4527), .A0(N18818), .A1(N4463), .B0(N2250), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3360 (.Y(N4528), .A0(N18818), .A1(N4464), .B0(N2251), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3361 (.Y(N4529), .A0(N18818), .A1(N4465), .B0(N2253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3362 (.Y(N4530), .A0(N18818), .A1(N4466), .B0(N2256), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3363 (.Y(N4531), .A0(N18818), .A1(N4467), .B0(N2257), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3364 (.Y(N4532), .A0(N18818), .A1(N4468), .B0(N2258), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3365 (.Y(N4533), .A0(N18818), .A1(N4469), .B0(N2259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I3366 (.Y(N4534), .A0(N18818), .A1(N4470), .B0(N2261), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I3367 (.Y(N4535), .A(inst_noninc_a_cellmath__55_2WWMM_in0[20]), .B(N4473));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4119 (.Y(N18331), .A0(N18544), .A1(N18227), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4121 (.Y(N5537), .A0(N18544), .A1(N18581), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4129 (.Y(N5550), .A0(N18544), .A1(N18219), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4131 (.Y(N18333), .A0(N18544), .A1(N18581), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4132 (.Y(N5553), .A0(N18544), .A1(N18405), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4133 (.Y(N5554), .A0(N18544), .A1(N18219), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4134 (.Y(N5555), .A(N18544), .B(N18589));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4135 (.Y(N5558), .A0(N18544), .A1(N18405), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4138 (.Y(N18335), .A0(N18544), .A1(N18589), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4139 (.Y(N18337), .A0(N18544), .A1(N18217), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4141 (.Y(N18339), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I4142 (.Y(N18341), .A(N18544), .B(N18416));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4150 (.Y(N5578), .A(N18544), .B(N18227));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4152 (.Y(N5584), .A0(N18544), .A1(N18581), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4153 (.Y(N18343), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4154 (.Y(N5586), .A0(N18544), .A1(N18589), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4157 (.Y(N5591), .A0(N18544), .A1(N18581), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4158 (.Y(N5592), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4159 (.Y(N5593), .A0(N18544), .A1(N18581), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I4160 (.Y(N5594), .A(N18223));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4161 (.Y(N18345), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4164 (.Y(N18347), .A0(N18544), .A1(N18424), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4933 (.Y(N6610), .A0(N18544), .A1(N18424), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4934 (.Y(N18349), .A0(N18544), .A1(N18424), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4936 (.Y(N6613), .A0(N18544), .A1(N18405), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I4949 (.Y(N6633), .A(N18544), .B(N18589));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I4950 (.Y(N6635), .A(N18581), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4952 (.Y(N6638), .A0(N18544), .A1(N18225), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4955 (.Y(N6641), .A0(N18544), .A1(N18225), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4956 (.Y(N6642), .A0(N18544), .A1(N18589), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4957 (.Y(N6643), .A0(N18544), .A1(N18416), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I4961 (.Y(N6648), .A(N18221));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4963 (.Y(N18351), .A(N18544), .B(inst_noninc_a_cellmath__55_2WWMM_in0[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4965 (.Y(N18353), .A0(N18544), .A1(N18405), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4966 (.Y(N6657), .A0(N18544), .A1(N18416), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4967 (.Y(N18355), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4975 (.Y(N6670), .A0(N18714), .A1(N18337), .B0(N18331), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4976 (.Y(N6671), .A0(N18714), .A1(N4351), .B0(N18259), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4977 (.Y(N6672), .A0(N18714), .A1(N18311), .B0(N5537), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4978 (.Y(N6673), .A0(N18714), .A1(N18343), .B0(N18313), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4985 (.Y(N6683), .A0(N18714), .A1(N18281), .B0(N5550), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4986 (.Y(N6684), .A0(N18714), .A1(N1103), .B0(N18325), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4987 (.Y(N6685), .A0(N18714), .A1(N6610), .B0(N18333), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4988 (.Y(N6686), .A0(N18714), .A1(N18349), .B0(N5553), .B1(N19053));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I4989 (.Y(N6687), .A(N18714), .B(N5554));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4990 (.Y(N6690), .A0(N18714), .A1(N6613), .B0(N5555), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4991 (.Y(N6691), .A0(N18714), .A1(N18239), .B0(N5558), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4992 (.Y(N6692), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18313), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4993 (.Y(N6693), .A0(N18714), .A1(N18557), .B0(N18277), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4994 (.Y(N6694), .A0(N18714), .A1(N18265), .B0(N18335), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4995 (.Y(N6695), .A0(N18714), .A1(N18311), .B0(N18337), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4996 (.Y(N6696), .A0(N18714), .A1(N18335), .B0(N18275), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4997 (.Y(N6697), .A0(N18714), .A1(N18315), .B0(N18339), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I4998 (.Y(N6698), .A0(N18714), .A1(N18267), .B0(N18341), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5003 (.Y(N6707), .A0(N18714), .A1(N6633), .B0(N18317), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5004 (.Y(N6708), .A0(N18714), .A1(N6635), .B0(N18301), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5005 (.Y(N6709), .A0(N18714), .A1(N18287), .B0(N18265), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5006 (.Y(N6710), .A0(N18714), .A1(N6638), .B0(N5578), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5007 (.Y(N6711), .A0(N18714), .A1(N18297), .B0(N18245), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5008 (.Y(N6712), .A0(N18714), .A1(N18333), .B0(N5584), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5009 (.Y(N6713), .A0(N18714), .A1(N6641), .B0(N18343), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5010 (.Y(N6714), .A0(N18714), .A1(N6642), .B0(N5586), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5011 (.Y(N6715), .A0(N18714), .A1(N6643), .B0(N2163), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5012 (.Y(N6716), .A0(N18714), .A1(N5591), .B0(N18341), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5013 (.Y(N6717), .A0(N18714), .A1(N18235), .B0(N5591), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5014 (.Y(N6718), .A0(N18714), .A1(N18341), .B0(N5592), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5015 (.Y(N6719), .A0(N18714), .A1(N6648), .B0(N5593), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5016 (.Y(N6720), .A0(N18714), .A1(N2163), .B0(N5594), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5017 (.Y(N6721), .A0(N18714), .A1(N18351), .B0(N18345), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5018 (.Y(N6722), .A0(N18714), .A1(N18257), .B0(N18279), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5019 (.Y(N6723), .A0(N18714), .A1(N18353), .B0(N18309), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5020 (.Y(N6724), .A0(N18714), .A1(N6657), .B0(N18347), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5021 (.Y(N6725), .A0(N18714), .A1(N18355), .B0(N18309), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5022 (.Y(N6726), .A0(N18714), .A1(N18313), .B0(N18271), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5023 (.Y(N6727), .A0(N18714), .A1(N18247), .B0(N18323), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I5778 (.Y(N7736), .A(N18219), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5779 (.Y(N18357), .A0(N18544), .A1(N18405), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5780 (.Y(N7739), .A0(N18544), .A1(N18589), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5787 (.Y(N7753), .A0(N18544), .A1(N18219), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I5789 (.Y(N7755), .A(N18581));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5793 (.Y(N7759), .A0(N18544), .A1(N18225), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5806 (.Y(N7780), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5808 (.Y(N7783), .A0(N18544), .A1(N18217), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5815 (.Y(N7790), .A0(N18544), .A1(N18416), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I5820 (.Y(N7795), .A(N18544), .B(N18215));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5823 (.Y(N7799), .A0(N18544), .A1(N18227), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6579 (.Y(N8814), .A0(N18544), .A1(N18227), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6581 (.Y(N18359), .A0(N18544), .A1(N18589), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6583 (.Y(N8819), .A0(N18544), .A1(N18221), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6590 (.Y(N8831), .A0(N18544), .A1(N18225), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6597 (.Y(N8843), .A0(N18544), .A1(N18223), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6599 (.Y(N8845), .A0(N18544), .A1(N18424), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6608 (.Y(N8861), .A0(N18544), .A1(N18217), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I6609 (.Y(N8862), .A(N18227));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6610 (.Y(N8863), .A(N18217), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6613 (.Y(N8867), .A0(N18544), .A1(N18225), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6614 (.Y(N8868), .A0(N18544), .A1(N18223), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6616 (.Y(N8870), .A0(N18544), .A1(N18217), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6617 (.Y(N8871), .A0(N18544), .A1(N18219), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6619 (.Y(N8873), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18405));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6624 (.Y(N18361), .A0(N18544), .A1(N18221), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6633 (.Y(N8895), .A0(N18714), .A1(N8814), .B0(N18327), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6634 (.Y(N8896), .A0(N18714), .A1(N18341), .B0(N7736), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6635 (.Y(N8897), .A0(N18714), .A1(N18359), .B0(N18357), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6636 (.Y(N8898), .A0(N18714), .A1(N18319), .B0(N7739), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6637 (.Y(N8899), .A0(N18714), .A1(N8819), .B0(N18301), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6638 (.Y(N8900), .A0(N18714), .A1(N18231), .B0(N18301), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6639 (.Y(N8901), .A(N18301), .B(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6643 (.Y(N8909), .A0(N18714), .A1(N6610), .B0(N7753), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6644 (.Y(N8910), .A0(N18714), .A1(N8831), .B0(N18337), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6645 (.Y(N8911), .A0(N18714), .A1(N5578), .B0(N7755), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6646 (.Y(N8912), .A0(N18714), .A1(N5558), .B0(N2180), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6647 (.Y(N8913), .A0(N18714), .A1(N5578), .B0(N18325), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6648 (.Y(N8914), .A0(N18714), .A1(N4371), .B0(N2179), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6649 (.Y(N8915), .A0(N18714), .A1(N2175), .B0(N7759), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6650 (.Y(N8916), .A0(N18714), .A1(N18279), .B0(N7736), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6651 (.Y(N8917), .A(N18714), .B(N8843));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6652 (.Y(N8919), .A(N19053), .B(N18255));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6653 (.Y(N8922), .A0(N18714), .A1(N8845), .B0(N18405), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6654 (.Y(N8923), .A0(N18714), .A1(N18319), .B0(N18607), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6655 (.Y(N8924), .A0(N18714), .A1(N18271), .B0(N18265), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6656 (.Y(N8925), .A0(N18714), .A1(N18247), .B0(N18269), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6657 (.Y(N8926), .A(N19055), .B(N18341));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6661 (.Y(N8933), .A0(N18714), .A1(N18327), .B0(N1068), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6662 (.Y(N8934), .A0(N18714), .A1(N8861), .B0(N7780), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6663 (.Y(N8935), .A0(N18714), .A1(N8862), .B0(N18544), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6664 (.Y(N8936), .A0(N18714), .A1(N8863), .B0(N7783), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6665 (.Y(N8937), .A0(N18714), .A1(N1086), .B0(N18321), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6666 (.Y(N8938), .A0(N18714), .A1(N18289), .B0(N6638), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6667 (.Y(N8939), .A0(N18714), .A1(N8867), .B0(N5592), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6668 (.Y(N8940), .A0(N18714), .A1(N8868), .B0(N18331), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6669 (.Y(N8941), .A0(N18714), .A1(N18353), .B0(N18275), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6670 (.Y(N8942), .A0(N18714), .A1(N8870), .B0(N18277), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6671 (.Y(N8943), .A0(N18714), .A1(N8871), .B0(N7790), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6672 (.Y(N8944), .A0(N18714), .A1(N18337), .B0(N18255), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6673 (.Y(N8945), .A0(N18714), .A1(N8873), .B0(N1066), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6674 (.Y(N8946), .A0(N18714), .A1(N18331), .B0(N18273), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6675 (.Y(N8947), .A0(N18714), .A1(N6635), .B0(N18297), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6676 (.Y(N8948), .A0(N18714), .A1(N18355), .B0(N7795), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6677 (.Y(N8949), .A0(N18714), .A1(N18347), .B0(N18291), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6678 (.Y(N8950), .A0(N18714), .A1(N18361), .B0(N18349), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6679 (.Y(N8951), .A0(N18714), .A1(N18353), .B0(N7799), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6680 (.Y(N8952), .A0(N18714), .A1(N7739), .B0(N18275), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6681 (.Y(N8953), .A0(N18714), .A1(N18301), .B0(N18253), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6682 (.Y(N8954), .A0(N18714), .A1(N18231), .B0(N18253), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6687 (.Y(N8962), .A0(N18818), .A1(N8895), .B0(N6670), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6688 (.Y(N8963), .A0(N18818), .A1(N8896), .B0(N6671), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6689 (.Y(N8964), .A0(N18818), .A1(N8897), .B0(N6672), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6690 (.Y(N8965), .A0(N18818), .A1(N8898), .B0(N6673), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6691 (.Y(N8966), .A0(N18818), .A1(N8899), .B0(N4469), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6692 (.Y(N8967), .A0(N18818), .A1(N8900), .B0(N4473), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6693 (.Y(N8968), .A(N18818), .B(N8901));
NOR2XL andori2bb1_A_I14502 (.Y(N19150), .A(N18714), .B(N18231));
NOR2XL andori2bb1_A_I14503 (.Y(N8972), .A(N19150), .B(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6697 (.Y(N8977), .A0(N18818), .A1(N8909), .B0(N6683), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6698 (.Y(N8978), .A0(N18818), .A1(N8910), .B0(N6684), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6699 (.Y(N8979), .A0(N18818), .A1(N8911), .B0(N6685), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6700 (.Y(N8980), .A0(N18818), .A1(N8912), .B0(N6686), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6701 (.Y(N8981), .A0(N18818), .A1(N8913), .B0(N6687), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6702 (.Y(N8982), .A0(N18818), .A1(N8914), .B0(N6690), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6703 (.Y(N8983), .A0(N18818), .A1(N8915), .B0(N6691), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6704 (.Y(N8984), .A0(N18818), .A1(N8916), .B0(N6692), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6705 (.Y(N8985), .A0(N18818), .A1(N8917), .B0(N6693), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6706 (.Y(N8986), .A0(N18818), .A1(N8919), .B0(N6694), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6707 (.Y(N8987), .A0(N18818), .A1(N8922), .B0(N6695), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6708 (.Y(N8988), .A0(N18818), .A1(N8923), .B0(N6696), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6709 (.Y(N8989), .A0(N18818), .A1(N8924), .B0(N6697), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6710 (.Y(N8990), .A0(N18818), .A1(N8925), .B0(N6698), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6711 (.Y(N8991), .A0(N18818), .A1(N8926), .B0(N2261), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6715 (.Y(N8998), .A0(N18818), .A1(N8933), .B0(N6707), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6716 (.Y(N8999), .A0(N18818), .A1(N8934), .B0(N6708), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6717 (.Y(N9000), .A0(N18818), .A1(N8935), .B0(N6709), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6718 (.Y(N9001), .A0(N18818), .A1(N8936), .B0(N6710), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6719 (.Y(N9002), .A0(N18818), .A1(N8937), .B0(N6711), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6720 (.Y(N9003), .A0(N18818), .A1(N8938), .B0(N6712), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6721 (.Y(N9004), .A0(N18818), .A1(N8939), .B0(N6713), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6722 (.Y(N9005), .A0(N18818), .A1(N8940), .B0(N6714), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6723 (.Y(N9006), .A0(N18818), .A1(N8941), .B0(N6715), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6724 (.Y(N9007), .A0(N18818), .A1(N8942), .B0(N6716), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6725 (.Y(N9008), .A0(N18818), .A1(N8943), .B0(N6717), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6726 (.Y(N9009), .A0(N18818), .A1(N8944), .B0(N6718), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6727 (.Y(N9010), .A0(N18818), .A1(N8945), .B0(N6719), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6728 (.Y(N9011), .A0(N18818), .A1(N8946), .B0(N6720), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6729 (.Y(N9012), .A0(N18818), .A1(N8947), .B0(N6721), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6730 (.Y(N9013), .A0(N18818), .A1(N8948), .B0(N6722), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6731 (.Y(N9014), .A0(N18818), .A1(N8949), .B0(N6723), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6732 (.Y(N9015), .A0(N18818), .A1(N8950), .B0(N6724), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6733 (.Y(N9016), .A0(N18818), .A1(N8951), .B0(N6725), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6734 (.Y(N9017), .A0(N18818), .A1(N8952), .B0(N6726), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6735 (.Y(N9018), .A0(N18818), .A1(N8953), .B0(N6727), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6736 (.Y(N9019), .A0(N18818), .A1(N8954), .B0(N19055), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I14485 (.Y(N9020), .A0N(N18253), .A1N(N19055), .B0(N18818));
NOR2XL andori2bb1_A_I14504 (.Y(N19157), .A(N18714), .B(N18323));
NOR2XL andori2bb1_A_I14505 (.Y(N9022), .A(N19157), .B(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I14210 (.Y(N18881), .A(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6741 (.Y(N9028), .A0(N18881), .A1(N8962), .B0(N4478), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6742 (.Y(N9029), .A0(N18881), .A1(N8963), .B0(N4479), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6743 (.Y(N9030), .A0(N18881), .A1(N8964), .B0(N4480), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6744 (.Y(N9031), .A0(N18881), .A1(N8965), .B0(N4481), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6745 (.Y(N9032), .A0(N18881), .A1(N8966), .B0(N4482), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6746 (.Y(N9033), .A0(N18881), .A1(N8967), .B0(N4483), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6747 (.Y(N9034), .A(N18881), .B(N8968));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I6748 (.Y(N9036), .A(inst_noninc_a_cellmath__55_2WWMM_in0[21]), .B(N8968));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6749 (.Y(N9039), .A(N18881), .B(N8972));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6751 (.Y(N9042), .A0(N18881), .A1(N8977), .B0(N4493), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6752 (.Y(N9043), .A0(N18881), .A1(N8978), .B0(N4494), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6753 (.Y(N9044), .A0(N18881), .A1(N8979), .B0(N4495), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6754 (.Y(N9045), .A0(N18881), .A1(N8980), .B0(N4496), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6755 (.Y(N9046), .A0(N18881), .A1(N8981), .B0(N4497), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6756 (.Y(N9047), .A0(N18881), .A1(N8982), .B0(N4498), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6757 (.Y(N9048), .A0(N18881), .A1(N8983), .B0(N4499), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6758 (.Y(N9049), .A0(N18881), .A1(N8984), .B0(N4500), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6759 (.Y(N9050), .A0(N18881), .A1(N8985), .B0(N4501), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6760 (.Y(N9051), .A0(N18881), .A1(N8986), .B0(N4502), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6761 (.Y(N9052), .A0(N18881), .A1(N8987), .B0(N4503), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6762 (.Y(N9053), .A0(N18881), .A1(N8988), .B0(N4504), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6763 (.Y(N9054), .A0(N18881), .A1(N8989), .B0(N4505), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6764 (.Y(N9055), .A0(N18881), .A1(N8990), .B0(N4506), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6765 (.Y(N9056), .A0(N18881), .A1(N8991), .B0(N4507), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
NOR2XL andori2bb1_A_I14506 (.Y(N19164), .A(N18818), .B(N18283));
NOR2XL andori2bb1_A_I14507 (.Y(N9057), .A(N19164), .B(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6769 (.Y(N9063), .A0(N18881), .A1(N8998), .B0(N4513), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6770 (.Y(N9064), .A0(N18881), .A1(N8999), .B0(N4514), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6771 (.Y(N9065), .A0(N18881), .A1(N9000), .B0(N4515), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6772 (.Y(N9066), .A0(N18881), .A1(N9001), .B0(N4516), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6773 (.Y(N9067), .A0(N18881), .A1(N9002), .B0(N4517), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6774 (.Y(N9068), .A0(N18881), .A1(N9003), .B0(N4518), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6775 (.Y(N9069), .A0(N18881), .A1(N9004), .B0(N4519), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6776 (.Y(N9070), .A0(N18881), .A1(N9005), .B0(N4520), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6777 (.Y(N9071), .A0(N18881), .A1(N9006), .B0(N4521), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6778 (.Y(N9072), .A0(N18881), .A1(N9007), .B0(N4522), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6779 (.Y(N9073), .A0(N18881), .A1(N9008), .B0(N4523), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6780 (.Y(N9074), .A0(N18881), .A1(N9009), .B0(N4524), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6781 (.Y(N9075), .A0(N18881), .A1(N9010), .B0(N4525), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6782 (.Y(N9076), .A0(N18881), .A1(N9011), .B0(N4526), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6783 (.Y(N9077), .A0(N18881), .A1(N9012), .B0(N4527), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6784 (.Y(N9078), .A0(N18881), .A1(N9013), .B0(N4528), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6785 (.Y(N9079), .A0(N18881), .A1(N9014), .B0(N4529), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6786 (.Y(N9080), .A0(N18881), .A1(N9015), .B0(N4530), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6787 (.Y(N9081), .A0(N18881), .A1(N9016), .B0(N4531), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6788 (.Y(N9082), .A0(N18881), .A1(N9017), .B0(N4532), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6789 (.Y(N9083), .A0(N18881), .A1(N9018), .B0(N4533), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6790 (.Y(N9084), .A0(N18881), .A1(N9019), .B0(N4534), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6791 (.Y(N9085), .A0(N18881), .A1(N9020), .B0(N4535), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I6792 (.Y(N9086), .A(N18881), .B(N9022));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7559 (.Y(N10112), .A0(N18544), .A1(N18405), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7575 (.Y(N10134), .A0(N18544), .A1(N18589), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7577 (.Y(N10137), .A0(N18544), .A1(N18223), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I7584 (.Y(N10146), .A0(N18544), .A1(N18215), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8348 (.Y(N11159), .A0(N18544), .A1(N18581), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8361 (.Y(N11176), .A(N18416), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I8362 (.Y(N11178), .A(N18544), .B(N18405));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8363 (.Y(N11181), .A(N18589), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8377 (.Y(N11204), .A0(N18544), .A1(N18215), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8379 (.Y(N11207), .A0(N18544), .A1(N18221), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8382 (.Y(N11210), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8399 (.Y(N11236), .A0(N18714), .A1(N18341), .B0(N7799), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8400 (.Y(N11237), .A0(N18714), .A1(N18359), .B0(N3314), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8401 (.Y(N11238), .A0(N18714), .A1(N18229), .B0(N18259), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8402 (.Y(N11239), .A0(N18714), .A1(N11159), .B0(N5537), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8403 (.Y(N11240), .A0(N18714), .A1(N7790), .B0(N18271), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8404 (.Y(N11241), .A0(N18714), .A1(N18239), .B0(N18253), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8405 (.Y(N11242), .A0(N18714), .A1(N18341), .B0(N18323), .B1(N19055));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8406 (.Y(N11243), .A(N18714), .B(N18247));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8409 (.Y(N11248), .A0(N18714), .A1(N1084), .B0(N18343), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8410 (.Y(N11249), .A0(N18714), .A1(N6641), .B0(N4342), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8411 (.Y(N11250), .A0(N18714), .A1(N18233), .B0(N18297), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8412 (.Y(N11251), .A0(N18714), .A1(N5558), .B0(N18357), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8413 (.Y(N11252), .A0(N18714), .A1(N4377), .B0(N4367), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8414 (.Y(N11253), .A0(N18714), .A1(N4377), .B0(N5554), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8415 (.Y(N11254), .A0(N18714), .A1(N11176), .B0(N10112), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8416 (.Y(N11255), .A0(N18714), .A1(N11178), .B0(N18341), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8417 (.Y(N11256), .A0(N18714), .A1(N11181), .B0(N18405), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8418 (.Y(N11257), .A0(N18714), .A1(N18357), .B0(N18607), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8419 (.Y(N11258), .A0(N18714), .A1(N18607), .B0(N18325), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8420 (.Y(N11259), .A0(N18714), .A1(N18321), .B0(N18279), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8427 (.Y(N11271), .A0(N18714), .A1(N8861), .B0(N18339), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8428 (.Y(N11272), .A0(N18714), .A1(N3314), .B0(N18291), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8429 (.Y(N11273), .A0(N18714), .A1(N18353), .B0(N18307), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8430 (.Y(N11274), .A0(N18714), .A1(N18247), .B0(N10112), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8431 (.Y(N11275), .A0(N18714), .A1(N11204), .B0(N10134), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8432 (.Y(N11276), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8433 (.Y(N11277), .A0(N18714), .A1(N11207), .B0(N10137), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8434 (.Y(N11278), .A0(N18714), .A1(N11207), .B0(N8862), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8435 (.Y(N11279), .A0(N18714), .A1(N18321), .B0(N3306), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8436 (.Y(N11280), .A0(N18714), .A1(N11210), .B0(N18273), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8437 (.Y(N11281), .A0(N18714), .A1(N18544), .B0(N18243), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8438 (.Y(N11282), .A0(N18714), .A1(N5550), .B0(N18309), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8439 (.Y(N11283), .A0(N18714), .A1(N18259), .B0(N18305), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8440 (.Y(N11284), .A0(N18714), .A1(N5553), .B0(N10146), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8441 (.Y(N11285), .A0(N18714), .A1(N2140), .B0(N18345), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8442 (.Y(N11286), .A0(N18714), .A1(N18267), .B0(N18279), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I8443 (.Y(N11287), .A(N18361), .B(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8445 (.Y(N11292), .A0(N18714), .A1(N18405), .B0(N18345), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8446 (.Y(N11293), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N7790), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8447 (.Y(N11294), .A0(N18714), .A1(N1102), .B0(N18239), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I8448 (.Y(N11295), .A0(N18714), .A1(N18247), .B0(N18341), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I8449 (.Y(N11296), .A(N18714), .B(N18247));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I9211 (.Y(N12316), .A(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9213 (.Y(N12319), .A0(N18544), .A1(N18227), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9218 (.Y(N12328), .A0(N18544), .A1(N18416), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I9229 (.Y(N12343), .A(N18544), .B(N18217));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9230 (.Y(N12346), .A0(N18544), .A1(N18221), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9237 (.Y(N12357), .A0(N18544), .A1(N18217), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9240 (.Y(N12362), .A0(N18544), .A1(N18217), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I9241 (.Y(N12363), .A(N18544), .B(N18223));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I9242 (.Y(N12366), .A0(N18544), .A1(N18215), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I9243 (.Y(N12367), .A(N18223), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10013 (.Y(N13404), .A(N18544), .B(N18223));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10014 (.Y(N13406), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10015 (.Y(N13407), .A0(N18544), .A1(N18227), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I10016 (.Y(N13408), .A(N18544), .B(N18424));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10017 (.Y(N13411), .A0(N18544), .A1(N18215), .B0(N18217), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10032 (.Y(N13437), .A0(N18544), .A1(N18416), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10036 (.Y(N13443), .A0(N18544), .A1(N18223), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10040 (.Y(N13448), .A0(N18544), .A1(N18217), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10048 (.Y(N13459), .A0(N18544), .A1(N18424), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10051 (.Y(N13462), .A0(N18544), .A1(N18215), .B0(N18219), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10057 (.Y(N13471), .A0(N18714), .A1(N1044), .B0(N4350), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10058 (.Y(N13472), .A0(N18714), .A1(N7739), .B0(N18351), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10059 (.Y(N13473), .A0(N18714), .A1(N18231), .B0(N18285), .B1(N19055));
INVXL inst_noninc_a_cellmath__55_2WWMM_I10061 (.Y(N13476), .A(N18557));
INVXL inst_noninc_a_cellmath__55_2WWMM_I10062 (.Y(N13477), .A(N18281));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10063 (.Y(N13478), .A0(N18714), .A1(N18269), .B0(N18267), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10067 (.Y(N13487), .A0(N18714), .A1(N13404), .B0(N12316), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10068 (.Y(N13488), .A0(N18714), .A1(N13406), .B0(N18299), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10069 (.Y(N13489), .A0(N18714), .A1(N13407), .B0(N12319), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10070 (.Y(N13490), .A0(N18714), .A1(N13408), .B0(N18347), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10071 (.Y(N13491), .A0(N18714), .A1(N13411), .B0(N18245), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10072 (.Y(N13492), .A0(N18714), .A1(N18331), .B0(N18351), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10073 (.Y(N13493), .A0(N18714), .A1(N18353), .B0(N4380), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10074 (.Y(N13494), .A0(N18714), .A1(N5554), .B0(N12328), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10075 (.Y(N13495), .A0(N18714), .A1(N12343), .B0(N18293), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10076 (.Y(N13496), .A0(N18714), .A1(N18253), .B0(N18295), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10077 (.Y(N13497), .A0(N18714), .A1(N18323), .B0(N4351), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10078 (.Y(N13498), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N6610), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10079 (.Y(N13499), .A0(N18714), .A1(N18416), .B0(N2180), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10081 (.Y(N13501), .A0(N18714), .A1(N18247), .B0(N18301), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10085 (.Y(N13508), .A0(N18714), .A1(N2142), .B0(N12343), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10086 (.Y(N13509), .A0(N18714), .A1(N13437), .B0(N12346), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10087 (.Y(N13510), .A0(N18714), .A1(N2147), .B0(N12343), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10088 (.Y(N13511), .A0(N18714), .A1(N18333), .B0(N18359), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10089 (.Y(N13512), .A0(N18714), .A1(N18253), .B0(N18345), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10090 (.Y(N13513), .A0(N18714), .A1(N13443), .B0(N18313), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10091 (.Y(N13514), .A0(N18714), .A1(N12367), .B0(N7783), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10092 (.Y(N13515), .A0(N18714), .A1(N7799), .B0(N3309), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10093 (.Y(N13516), .A0(N18714), .A1(N1084), .B0(N12357), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10094 (.Y(N13517), .A0(N18714), .A1(N13448), .B0(N3306), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10095 (.Y(N13518), .A0(N18714), .A1(N18339), .B0(N18361), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10096 (.Y(N13519), .A0(N18714), .A1(N18239), .B0(N12362), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10097 (.Y(N13520), .A0(N18714), .A1(N18557), .B0(N12363), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10098 (.Y(N13521), .A0(N18714), .A1(N6642), .B0(N12366), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10099 (.Y(N13522), .A0(N18714), .A1(N18351), .B0(N12367), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10100 (.Y(N13523), .A0(N18714), .A1(N12367), .B0(N18345), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10101 (.Y(N13524), .A0(N18714), .A1(N18353), .B0(N18343), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10102 (.Y(N13525), .A0(N18714), .A1(N13459), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10103 (.Y(N13526), .A0(N18714), .A1(N18325), .B0(N4329), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10104 (.Y(N13527), .A0(N18714), .A1(N18305), .B0(N18293), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10105 (.Y(N13528), .A0(N18714), .A1(N13462), .B0(N18361), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10106 (.Y(N13529), .A0(N18714), .A1(N18544), .B0(N18301), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10111 (.Y(N13538), .A0(N18818), .A1(N13471), .B0(N11236), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10112 (.Y(N13539), .A0(N18818), .A1(N13472), .B0(N11237), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10113 (.Y(N13540), .A0(N18818), .A1(N13473), .B0(N11238), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10114 (.Y(N13541), .A0(N18818), .A1(N18405), .B0(N11239), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10115 (.Y(N13542), .A0(N18818), .A1(N13476), .B0(N11240), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10116 (.Y(N13543), .A0(N18818), .A1(N13477), .B0(N11241), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10117 (.Y(N13544), .A0(N18818), .A1(N13478), .B0(N11242), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10118 (.Y(N13545), .A0(N18818), .A1(N18283), .B0(N11243), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10119 (.Y(N13546), .A(N18818), .B(N18283));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10121 (.Y(N13551), .A0(N18818), .A1(N13487), .B0(N11248), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10122 (.Y(N13552), .A0(N18818), .A1(N13488), .B0(N11249), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10123 (.Y(N13553), .A0(N18818), .A1(N13489), .B0(N11250), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10124 (.Y(N13554), .A0(N18818), .A1(N13490), .B0(N11251), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10125 (.Y(N13555), .A0(N18818), .A1(N13491), .B0(N11252), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10126 (.Y(N13556), .A0(N18818), .A1(N13492), .B0(N11253), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10127 (.Y(N13557), .A0(N18818), .A1(N13493), .B0(N11254), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10128 (.Y(N13558), .A0(N18818), .A1(N13494), .B0(N11255), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10129 (.Y(N13559), .A0(N18818), .A1(N13495), .B0(N11256), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10130 (.Y(N13560), .A0(N18818), .A1(N13496), .B0(N11257), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10131 (.Y(N13561), .A0(N18818), .A1(N13497), .B0(N11258), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10132 (.Y(N13562), .A0(N18818), .A1(N13498), .B0(N11259), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10133 (.Y(N13563), .A0(N18818), .A1(N13499), .B0(N4436), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10134 (.Y(N13564), .A0(N18818), .A1(N2202), .B0(N4437), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10135 (.Y(N13565), .A0(N18818), .A1(N13501), .B0(N18329), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10136 (.Y(N13566), .A0(N18818), .A1(N8926), .B0(N18329), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I10137 (.Y(N13567), .A(N18329), .B(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I10138 (.Y(N13569), .A(N18818), .B(N2253));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10139 (.Y(N13572), .A0(N18818), .A1(N13508), .B0(N11271), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10140 (.Y(N13573), .A0(N18818), .A1(N13509), .B0(N11272), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10141 (.Y(N13574), .A0(N18818), .A1(N13510), .B0(N11273), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10142 (.Y(N13575), .A0(N18818), .A1(N13511), .B0(N11274), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10143 (.Y(N13576), .A0(N18818), .A1(N13512), .B0(N11275), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10144 (.Y(N13577), .A0(N18818), .A1(N13513), .B0(N11276), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10145 (.Y(N13578), .A0(N18818), .A1(N13514), .B0(N11277), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10146 (.Y(N13579), .A0(N18818), .A1(N13515), .B0(N11278), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10147 (.Y(N13580), .A0(N18818), .A1(N13516), .B0(N11279), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10148 (.Y(N13581), .A0(N18818), .A1(N13517), .B0(N11280), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10149 (.Y(N13582), .A0(N18818), .A1(N13518), .B0(N11281), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10150 (.Y(N13583), .A0(N18818), .A1(N13519), .B0(N11282), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10151 (.Y(N13584), .A0(N18818), .A1(N13520), .B0(N11283), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10152 (.Y(N13585), .A0(N18818), .A1(N13521), .B0(N11284), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10153 (.Y(N13586), .A0(N18818), .A1(N13522), .B0(N11285), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10154 (.Y(N13587), .A0(N18818), .A1(N13523), .B0(N11286), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10155 (.Y(N13588), .A0(N18818), .A1(N13524), .B0(N11287), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10156 (.Y(N13589), .A0(N18818), .A1(N13525), .B0(N4417), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10157 (.Y(N13590), .A0(N18818), .A1(N13526), .B0(N11292), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10158 (.Y(N13591), .A0(N18818), .A1(N13527), .B0(N11293), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10159 (.Y(N13592), .A0(N18818), .A1(N13528), .B0(N11294), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10160 (.Y(N13593), .A0(N18818), .A1(N13529), .B0(N11295), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10161 (.Y(N13594), .A0(N18818), .A1(N8901), .B0(N11296), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I10923 (.Y(N14617), .A(N18219));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10925 (.Y(N14619), .A0(N18544), .A1(N18219), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10927 (.Y(N14621), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10941 (.Y(N14638), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10944 (.Y(N14641), .A0(N18544), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10950 (.Y(N14649), .A0(N18544), .A1(N18217), .B0(N18581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I10956 (.Y(N14658), .A0(N18544), .A1(N18405), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11728 (.Y(N15695), .A0(N18544), .A1(N18227), .B0(N18225), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11738 (.Y(N15708), .A0(N18544), .A1(N18225), .B0(N18221), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11750 (.Y(N15724), .A0(N18544), .A1(N18223), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11751 (.Y(N15725), .A0(N18544), .A1(N18221), .B0(N18227), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11769 (.Y(N15750), .A0(N18714), .A1(N18289), .B0(N8868), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11770 (.Y(N15751), .A0(N18714), .A1(N5592), .B0(N6657), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11771 (.Y(N15752), .A0(N18714), .A1(N18303), .B0(N18355), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11772 (.Y(N15753), .A0(N18714), .A1(N7759), .B0(N18259), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11773 (.Y(N15754), .A0(N18714), .A1(N18277), .B0(N18289), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11774 (.Y(N15755), .A0(N18714), .A1(N18349), .B0(N18361), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11775 (.Y(N15756), .A0(N18714), .A1(N18315), .B0(N18231), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11779 (.Y(N15762), .A0(N18714), .A1(N4342), .B0(N14617), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11780 (.Y(N15763), .A0(N18714), .A1(N18259), .B0(N18287), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11781 (.Y(N15764), .A0(N18714), .A1(N4344), .B0(N14619), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11782 (.Y(N15765), .A0(N18714), .A1(N15695), .B0(N8819), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11783 (.Y(N15766), .A0(N18714), .A1(N18335), .B0(N14621), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11784 (.Y(N15767), .A0(N18714), .A1(N4344), .B0(N8867), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11785 (.Y(N15768), .A0(N18714), .A1(N18309), .B0(N13448), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11786 (.Y(N15769), .A0(N18714), .A1(N8873), .B0(N2175), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11787 (.Y(N15770), .A0(N18714), .A1(N4371), .B0(N18279), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11788 (.Y(N15771), .A0(N18714), .A1(N8845), .B0(N8843), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11789 (.Y(N15772), .A0(N18714), .A1(N18319), .B0(N18255), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11790 (.Y(N15773), .A0(N18714), .A1(N18259), .B0(N18359), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11791 (.Y(N15774), .A0(N18714), .A1(N18309), .B0(N8861), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11792 (.Y(N15775), .A0(N18714), .A1(N15708), .B0(N18255), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11793 (.Y(N15776), .A0(N18714), .A1(N18544), .B0(N18341), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11797 (.Y(N15783), .A0(N18714), .A1(N8845), .B0(N14638), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11798 (.Y(N15784), .A0(N18714), .A1(N18339), .B0(N18261), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11799 (.Y(N15785), .A0(N18714), .A1(N8831), .B0(N18339), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11800 (.Y(N15786), .A0(N18714), .A1(N18309), .B0(N14641), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11801 (.Y(N15787), .A0(N18714), .A1(N18355), .B0(N5555), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11802 (.Y(N15788), .A0(N18714), .A1(N15708), .B0(N18277), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11803 (.Y(N15789), .A0(N18714), .A1(N18325), .B0(N18333), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11804 (.Y(N15790), .A0(N18714), .A1(N15724), .B0(N18349), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11805 (.Y(N15791), .A0(N18714), .A1(N15725), .B0(N18235), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11806 (.Y(N15792), .A0(N18714), .A1(N15724), .B0(N14649), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11807 (.Y(N15793), .A0(N18714), .A1(N18357), .B0(N18311), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11808 (.Y(N15794), .A0(N18714), .A1(N11207), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11809 (.Y(N15795), .A0(N18714), .A1(N8863), .B0(N18261), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11810 (.Y(N15796), .A0(N18714), .A1(N18317), .B0(N1044), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11811 (.Y(N15797), .A0(N18714), .A1(N14649), .B0(N11176), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11812 (.Y(N15798), .A0(N18714), .A1(N8867), .B0(N14658), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11813 (.Y(N15799), .A0(N18714), .A1(N11204), .B0(N4396), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11814 (.Y(N15800), .A0(N18714), .A1(N18405), .B0(N18259), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11815 (.Y(N15801), .A0(N18714), .A1(N18557), .B0(N18305), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11816 (.Y(N15802), .A0(N18714), .A1(N18331), .B0(N18259), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11818 (.Y(N15804), .A0(N18714), .A1(N18341), .B0(N18285), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I11819 (.Y(N15805), .A0(N18714), .A1(N18341), .B0(N18257), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I12582 (.Y(N16832), .A(N18221), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12589 (.Y(N16845), .A0(N18544), .A1(N18227), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12601 (.Y(N16861), .A0(N18544), .A1(N18581), .B0(N18215), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12602 (.Y(N16862), .A0(N18544), .A1(N18217), .B0(N18405), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I12608 (.Y(N16869), .A(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B(N18581));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12612 (.Y(N16878), .A0(N18544), .A1(N18215), .B0(N18589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I12613 (.Y(N16879), .A(N18544), .B(N18424));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I12615 (.Y(N16882), .A0(N18544), .A1(N18405), .B0(N18416), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I13383 (.Y(N17901), .A(N18225));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13390 (.Y(N17908), .A(N18424), .B(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13413 (.Y(N17948), .A0(N18544), .A1(N18221), .B0(N18223), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13416 (.Y(N17951), .A0(N18544), .A1(N18221), .B0(N18424), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[18]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13427 (.Y(N17969), .A0(N18714), .A1(N5555), .B0(N18241), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13428 (.Y(N17970), .A0(N18714), .A1(N18317), .B0(N14658), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13429 (.Y(N17971), .A0(N18714), .A1(N18307), .B0(N6633), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13430 (.Y(N17972), .A0(N18714), .A1(N18305), .B0(N18231), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13431 (.Y(N17973), .A0(N18714), .A1(N18289), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[16]), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13432 (.Y(N17974), .A0(N18714), .A1(N18259), .B0(N18557), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13433 (.Y(N17975), .A0(N18714), .A1(N18299), .B0(N18265), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13434 (.Y(N17976), .A0(N18714), .A1(N18257), .B0(N18253), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13437 (.Y(N17982), .A0(N18714), .A1(N17901), .B0(N5593), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13438 (.Y(N17983), .A0(N18714), .A1(N18289), .B0(N16832), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13439 (.Y(N17984), .A0(N18714), .A1(N2141), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13440 (.Y(N17985), .A0(N18714), .A1(N16861), .B0(N12316), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13441 (.Y(N17986), .A0(N18714), .A1(N14619), .B0(N18243), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13442 (.Y(N17987), .A(N18714), .B(N10146));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13443 (.Y(N17989), .A0(N18714), .A1(N8814), .B0(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13444 (.Y(N17990), .A0(N18714), .A1(N17908), .B0(N2176), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13445 (.Y(N17991), .A0(N18714), .A1(N1089), .B0(N16845), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13446 (.Y(N17992), .A0(N18714), .A1(N18307), .B0(N18229), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13447 (.Y(N17993), .A0(N18714), .A1(N11181), .B0(N18333), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13448 (.Y(N17994), .A0(N18714), .A1(N1068), .B0(N18416), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13449 (.Y(N17995), .A0(N18714), .A1(N18357), .B0(N18291), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13450 (.Y(N17996), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[17]), .B0(N18335), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13451 (.Y(N17997), .A0(N18714), .A1(inst_noninc_a_cellmath__55_2WWMM_in0[18]), .B0(N18315), .B1(N19053));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13452 (.Y(N17998), .A(N18269), .B(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13455 (.Y(N18002), .A0(N18714), .A1(N18347), .B0(N14638), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13456 (.Y(N18003), .A0(N18714), .A1(N12363), .B0(N18271), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13457 (.Y(N18004), .A0(N18714), .A1(N1093), .B0(N16861), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13458 (.Y(N18005), .A0(N18714), .A1(N10134), .B0(N16862), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13459 (.Y(N18006), .A0(N18714), .A1(N7753), .B0(N4329), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13460 (.Y(N18007), .A0(N18714), .A1(N16878), .B0(N14649), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13461 (.Y(N18008), .A0(N18714), .A1(N18303), .B0(N18295), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13462 (.Y(N18009), .A0(N18714), .A1(N15724), .B0(N18301), .B1(N19053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13463 (.Y(N18010), .A0(N18714), .A1(N11210), .B0(N8819), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13464 (.Y(N18011), .A0(N18714), .A1(N11176), .B0(N16869), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13465 (.Y(N18012), .A0(N18714), .A1(N3309), .B0(N4382), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13466 (.Y(N18013), .A0(N18714), .A1(N1045), .B0(N18261), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13467 (.Y(N18014), .A0(N18714), .A1(N17948), .B0(N18245), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13468 (.Y(N18015), .A0(N18714), .A1(N18281), .B0(N16878), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13469 (.Y(N18016), .A0(N18714), .A1(N18295), .B0(N16879), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13470 (.Y(N18017), .A0(N18714), .A1(N17951), .B0(N12346), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13471 (.Y(N18018), .A0(N18714), .A1(N12363), .B0(N16882), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13472 (.Y(N18019), .A0(N18714), .A1(N18285), .B0(N3327), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13473 (.Y(N18020), .A(N18714), .B(N18327));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13474 (.Y(N18023), .A0(N18714), .A1(N18405), .B0(N18357), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13475 (.Y(N18024), .A0(N18714), .A1(N18416), .B0(N13459), .B1(N19055));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13476 (.Y(N18025), .A0(N18714), .A1(N18544), .B0(N18281), .B1(N19055));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13477 (.Y(N18026), .A(N18714), .B(N18267));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13481 (.Y(N18034), .A0(N18818), .A1(N17969), .B0(N15750), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13482 (.Y(N18035), .A0(N18818), .A1(N17970), .B0(N15751), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13483 (.Y(N18036), .A0(N18818), .A1(N17971), .B0(N15752), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13484 (.Y(N18037), .A0(N18818), .A1(N17972), .B0(N15753), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13485 (.Y(N18038), .A0(N18818), .A1(N17973), .B0(N15754), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13486 (.Y(N18039), .A0(N18818), .A1(N17974), .B0(N15755), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13487 (.Y(N18040), .A0(N18818), .A1(N17975), .B0(N15756), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13488 (.Y(N18041), .A0(N18818), .A1(N17976), .B0(N2203), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13491 (.Y(N18046), .A0(N18818), .A1(N17982), .B0(N15762), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13492 (.Y(N18047), .A0(N18818), .A1(N17983), .B0(N15763), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13493 (.Y(N18048), .A0(N18818), .A1(N17984), .B0(N15764), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13494 (.Y(N18049), .A0(N18818), .A1(N17985), .B0(N15765), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13495 (.Y(N18050), .A0(N18818), .A1(N17986), .B0(N15766), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13496 (.Y(N18051), .A0(N18818), .A1(N17987), .B0(N15767), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13497 (.Y(N18052), .A0(N18818), .A1(N17989), .B0(N15768), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13498 (.Y(N18053), .A0(N18818), .A1(N17990), .B0(N15769), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13499 (.Y(N18054), .A0(N18818), .A1(N17991), .B0(N15770), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13500 (.Y(N18055), .A0(N18818), .A1(N17992), .B0(N15771), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13501 (.Y(N18056), .A0(N18818), .A1(N17993), .B0(N15772), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13502 (.Y(N18057), .A0(N18818), .A1(N17994), .B0(N15773), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13503 (.Y(N18058), .A0(N18818), .A1(N17995), .B0(N15774), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13504 (.Y(N18059), .A0(N18818), .A1(N17996), .B0(N15775), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13505 (.Y(N18060), .A0(N18818), .A1(N17997), .B0(N15776), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13506 (.Y(N18061), .A0(N18818), .A1(N17998), .B0(N4473), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13507 (.Y(N18062), .A(N18818), .B(N4470));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13509 (.Y(N18067), .A0(N18818), .A1(N18002), .B0(N15783), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13510 (.Y(N18068), .A0(N18818), .A1(N18003), .B0(N15784), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13511 (.Y(N18069), .A0(N18818), .A1(N18004), .B0(N15785), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13512 (.Y(N18070), .A0(N18818), .A1(N18005), .B0(N15786), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13513 (.Y(N18071), .A0(N18818), .A1(N18006), .B0(N15787), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13514 (.Y(N18072), .A0(N18818), .A1(N18007), .B0(N15788), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13515 (.Y(N18073), .A0(N18818), .A1(N18008), .B0(N15789), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13516 (.Y(N18074), .A0(N18818), .A1(N18009), .B0(N15790), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13517 (.Y(N18075), .A0(N18818), .A1(N18010), .B0(N15791), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13518 (.Y(N18076), .A0(N18818), .A1(N18011), .B0(N15792), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13519 (.Y(N18077), .A0(N18818), .A1(N18012), .B0(N15793), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13520 (.Y(N18078), .A0(N18818), .A1(N18013), .B0(N15794), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13521 (.Y(N18079), .A0(N18818), .A1(N18014), .B0(N15795), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13522 (.Y(N18080), .A0(N18818), .A1(N18015), .B0(N15796), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13523 (.Y(N18081), .A0(N18818), .A1(N18016), .B0(N15797), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13524 (.Y(N18082), .A0(N18818), .A1(N18017), .B0(N15798), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13525 (.Y(N18083), .A0(N18818), .A1(N18018), .B0(N15799), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13526 (.Y(N18084), .A0(N18818), .A1(N18019), .B0(N15800), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13527 (.Y(N18085), .A0(N18818), .A1(N18020), .B0(N15801), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13528 (.Y(N18086), .A0(N18818), .A1(N18023), .B0(N15802), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13529 (.Y(N18087), .A0(N18818), .A1(N18024), .B0(N4436), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13530 (.Y(N18088), .A0(N18818), .A1(N18025), .B0(N15804), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13531 (.Y(N18089), .A0(N18818), .A1(N18026), .B0(N15805), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I13532 (.Y(N18090), .A(N11243), .B(inst_noninc_a_cellmath__55_2WWMM_in0[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13535 (.Y(N18094), .A0(N18881), .A1(N18034), .B0(N13538), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13536 (.Y(N18095), .A0(N18881), .A1(N18035), .B0(N13539), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13537 (.Y(N18096), .A0(N18881), .A1(N18036), .B0(N13540), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13538 (.Y(N18097), .A0(N18881), .A1(N18037), .B0(N13541), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13539 (.Y(N18098), .A0(N18881), .A1(N18038), .B0(N13542), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13540 (.Y(N18099), .A0(N18881), .A1(N18039), .B0(N13543), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13541 (.Y(N18100), .A0(N18881), .A1(N18040), .B0(N13544), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13542 (.Y(N18101), .A0(N18881), .A1(N18041), .B0(N13545), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13543 (.Y(N18102), .A0(N18881), .A1(N9022), .B0(N13546), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
NOR2XL andori2bb1_A_I14508 (.Y(N19171), .A(inst_noninc_a_cellmath__55_2WWMM_in0[20]), .B(N2261));
NOR2XL andori2bb1_A_I14509 (.Y(N18103), .A(N19171), .B(N18881));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13545 (.Y(N18106), .A0(N18881), .A1(N18046), .B0(N13551), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13546 (.Y(N18107), .A0(N18881), .A1(N18047), .B0(N13552), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13547 (.Y(N18108), .A0(N18881), .A1(N18048), .B0(N13553), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13548 (.Y(N18109), .A0(N18881), .A1(N18049), .B0(N13554), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13549 (.Y(N18110), .A0(N18881), .A1(N18050), .B0(N13555), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13550 (.Y(N18111), .A0(N18881), .A1(N18051), .B0(N13556), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13551 (.Y(N18112), .A0(N18881), .A1(N18052), .B0(N13557), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13552 (.Y(N18113), .A0(N18881), .A1(N18053), .B0(N13558), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13553 (.Y(N18114), .A0(N18881), .A1(N18054), .B0(N13559), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13554 (.Y(N18115), .A0(N18881), .A1(N18055), .B0(N13560), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13555 (.Y(N18116), .A0(N18881), .A1(N18056), .B0(N13561), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13556 (.Y(N18117), .A0(N18881), .A1(N18057), .B0(N13562), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13557 (.Y(N18118), .A0(N18881), .A1(N18058), .B0(N13563), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13558 (.Y(N18119), .A0(N18881), .A1(N18059), .B0(N13564), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13559 (.Y(N18120), .A0(N18881), .A1(N18060), .B0(N13565), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13560 (.Y(N18121), .A0(N18881), .A1(N18061), .B0(N13566), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13561 (.Y(N18122), .A0(N18881), .A1(N18062), .B0(N13567), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13563 (.Y(N18125), .A0(N18881), .A1(N18067), .B0(N13572), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13564 (.Y(N18126), .A0(N18881), .A1(N18068), .B0(N13573), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13565 (.Y(N18127), .A0(N18881), .A1(N18069), .B0(N13574), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13566 (.Y(N18128), .A0(N18881), .A1(N18070), .B0(N13575), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13567 (.Y(N18129), .A0(N18881), .A1(N18071), .B0(N13576), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13568 (.Y(N18130), .A0(N18881), .A1(N18072), .B0(N13577), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13569 (.Y(N18131), .A0(N18881), .A1(N18073), .B0(N13578), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13570 (.Y(N18132), .A0(N18881), .A1(N18074), .B0(N13579), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13571 (.Y(N18133), .A0(N18881), .A1(N18075), .B0(N13580), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13572 (.Y(N18134), .A0(N18881), .A1(N18076), .B0(N13581), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13573 (.Y(N18135), .A0(N18881), .A1(N18077), .B0(N13582), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13574 (.Y(N18136), .A0(N18881), .A1(N18078), .B0(N13583), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13575 (.Y(N18137), .A0(N18881), .A1(N18079), .B0(N13584), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13576 (.Y(N18138), .A0(N18881), .A1(N18080), .B0(N13585), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13577 (.Y(N18139), .A0(N18881), .A1(N18081), .B0(N13586), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13578 (.Y(N18140), .A0(N18881), .A1(N18082), .B0(N13587), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13579 (.Y(N18141), .A0(N18881), .A1(N18083), .B0(N13588), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13580 (.Y(N18142), .A0(N18881), .A1(N18084), .B0(N13589), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13581 (.Y(N18143), .A0(N18881), .A1(N18085), .B0(N13590), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13582 (.Y(N18144), .A0(N18881), .A1(N18086), .B0(N13591), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13583 (.Y(N18145), .A0(N18881), .A1(N18087), .B0(N13592), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13584 (.Y(N18146), .A0(N18881), .A1(N18088), .B0(N13593), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13585 (.Y(N18147), .A0(N18881), .A1(N18089), .B0(N13594), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13586 (.Y(N18148), .A0(N18881), .A1(N18090), .B0(N8968), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[21]));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I14225 (.Y(N18896), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13589 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[0]), .A0(N18896), .A1(N18094), .B0(N9028), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13590 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[1]), .A0(N18896), .A1(N18095), .B0(N9029), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13591 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[2]), .A0(N18896), .A1(N18096), .B0(N9030), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13592 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[3]), .A0(N18896), .A1(N18097), .B0(N9031), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13593 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[4]), .A0(N18896), .A1(N18098), .B0(N9032), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13594 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[5]), .A0(N18896), .A1(N18099), .B0(N9033), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13595 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[6]), .A0(N18896), .A1(N18100), .B0(N9034), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13596 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[7]), .A0(N18896), .A1(N18101), .B0(N9036), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13597 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[8]), .A0(N18896), .A1(N18102), .B0(N9039), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13598 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[9]), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]), .B(N18103));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13599 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[10]), .A0(N18896), .A1(N18106), .B0(N9042), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13600 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[11]), .A0(N18896), .A1(N18107), .B0(N9043), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13601 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[12]), .A0(N18896), .A1(N18108), .B0(N9044), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13602 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[13]), .A0(N18896), .A1(N18109), .B0(N9045), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13603 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[14]), .A0(N18896), .A1(N18110), .B0(N9046), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13604 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[15]), .A0(N18896), .A1(N18111), .B0(N9047), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13605 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[16]), .A0(N18896), .A1(N18112), .B0(N9048), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13606 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[17]), .A0(N18896), .A1(N18113), .B0(N9049), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13607 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[18]), .A0(N18896), .A1(N18114), .B0(N9050), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13608 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[19]), .A0(N18896), .A1(N18115), .B0(N9051), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13609 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[20]), .A0(N18896), .A1(N18116), .B0(N9052), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13610 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[21]), .A0(N18896), .A1(N18117), .B0(N9053), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13611 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[22]), .A0(N18896), .A1(N18118), .B0(N9054), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13612 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[23]), .A0(N18896), .A1(N18119), .B0(N9055), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13613 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[24]), .A0(N18896), .A1(N18120), .B0(N9056), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13614 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[25]), .A0(N18896), .A1(N18121), .B0(N9057), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I13615 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[26]), .A(inst_noninc_a_cellmath__55_2WWMM_in0[22]), .B(N18122));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I14489 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[27]), .A0N(N13569), .A1N(inst_noninc_a_cellmath__55_2WWMM_in0[21]), .B0(N18896));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13617 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[28]), .A0(N18896), .A1(N18125), .B0(N9063), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13618 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[29]), .A0(N18896), .A1(N18126), .B0(N9064), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13619 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[30]), .A0(N18896), .A1(N18127), .B0(N9065), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13620 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[31]), .A0(N18896), .A1(N18128), .B0(N9066), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13621 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[32]), .A0(N18896), .A1(N18129), .B0(N9067), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13622 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[33]), .A0(N18896), .A1(N18130), .B0(N9068), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13623 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[34]), .A0(N18896), .A1(N18131), .B0(N9069), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13624 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[35]), .A0(N18896), .A1(N18132), .B0(N9070), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13625 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[36]), .A0(N18896), .A1(N18133), .B0(N9071), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13626 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[37]), .A0(N18896), .A1(N18134), .B0(N9072), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13627 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[38]), .A0(N18896), .A1(N18135), .B0(N9073), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13628 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[39]), .A0(N18896), .A1(N18136), .B0(N9074), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13629 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[40]), .A0(N18896), .A1(N18137), .B0(N9075), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13630 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[41]), .A0(N18896), .A1(N18138), .B0(N9076), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13631 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[42]), .A0(N18896), .A1(N18139), .B0(N9077), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13632 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[43]), .A0(N18896), .A1(N18140), .B0(N9078), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13633 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[44]), .A0(N18896), .A1(N18141), .B0(N9079), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13634 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[45]), .A0(N18896), .A1(N18142), .B0(N9080), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13635 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[46]), .A0(N18896), .A1(N18143), .B0(N9081), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13636 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[47]), .A0(N18896), .A1(N18144), .B0(N9082), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13637 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[48]), .A0(N18896), .A1(N18145), .B0(N9083), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13638 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[49]), .A0(N18896), .A1(N18146), .B0(N9084), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13639 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[50]), .A0(N18896), .A1(N18147), .B0(N9085), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I13640 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[51]), .A0(N18896), .A1(N18148), .B0(N9086), .B1(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
NOR2XL andori2bb1_A_I14510 (.Y(N19178), .A(N18881), .B(N8972));
NOR2XL andori2bb1_A_I14511 (.Y(inst_noninc_a_cellmath__55_2WWMM_out0[52]), .A(N19178), .B(inst_noninc_a_cellmath__55_2WWMM_in0[22]));
endmodule

module cynw_cm_float_rcp_inst_cellmath__62_0_bdw1412651405_bdw (
	inst_cellmath__62_0_out0,
	inst_cellmath__62_0_out1,
	inst_cellmath__62_0_in0,
	inst_cellmath__62_0_in1
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__62_0_out0,
	inst_cellmath__62_0_out1;
input [9:0] inst_cellmath__62_0_in0;
input [24:13] inst_cellmath__62_0_in1;
wire N313,N315,N317,N319,N321,N323,N325 
	,N327,N329,N331,N348,N350,N352,N354,N356 
	,N358,N360,N362,N364,N366,N379,N381,N383 
	,N385,N387,N389,N391,N393,N395,N397,N399 
	,N401,N414,N416,N418,N420,N422,N424,N426 
	,N428,N430,N432,N434,N436,N449,N451,N453 
	,N455,N457,N459,N461,N463,N465,N467,N469 
	,N471,N484,N486,N488,N490,N492,N494,N496 
	,N498,N500,N502,N504,N506,N519,N521,N523 
	,N525,N527,N529,N531,N533,N535,N537,N539 
	,N541,N554,N556,N558,N560,N562,N564,N566 
	,N568,N570,N572,N574,N576,N589,N591,N593 
	,N595,N597,N599,N601,N603,N605,N607,N609 
	,N611,N624,N626,N628,N630,N632,N634,N636 
	,N638,N640,N642,N644,N650,N652,N654,N655 
	,N656,N658,N661,N662,N663,N664,N665,N666 
	,N669,N670,N671,N672,N673,N674,N675,N676 
	,N679,N680,N681,N682,N683,N684,N685,N686 
	,N687,N688,N691,N692,N693,N694,N695,N696 
	,N697,N698,N699,N700,N701,N702,N705,N706 
	,N707,N708,N709,N710,N711,N712,N713,N714 
	,N715,N716,N717,N718,N721,N722,N723,N724 
	,N725,N726,N727,N728,N729,N730,N731,N732 
	,N733,N734,N737,N738,N739,N740,N741,N742 
	,N743,N744,N745,N746,N747,N748,N749,N750 
	,N753,N754,N755,N756,N757,N758,N759,N760 
	,N761,N762,N763,N764,N765,N766,N769,N770 
	,N771,N772,N773,N774,N775,N776,N777,N778 
	,N779,N780,N783,N784,N785,N786,N787,N788 
	,N789,N790,N791,N792,N795,N796,N797,N798 
	,N799,N800,N801,N802,N805,N806,N807,N808 
	,N809,N810,N813,N814,N815,N816,N819,N820 
	,N825,N826,N827,N828,N829,N830,N831,N832 
	,N833,N834,N835,N836,N837,N838,N839,N840 
	,N841,N842,N843,N844,N845,N846;
INVXL inst_cellmath__62_0_I303 (.Y(N825), .A(inst_cellmath__62_0_in1[13]));
INVXL inst_cellmath__62_0_I304 (.Y(N826), .A(inst_cellmath__62_0_in1[14]));
INVXL inst_cellmath__62_0_I305 (.Y(N827), .A(inst_cellmath__62_0_in1[15]));
INVXL inst_cellmath__62_0_I306 (.Y(N828), .A(inst_cellmath__62_0_in1[16]));
INVXL inst_cellmath__62_0_I307 (.Y(N829), .A(inst_cellmath__62_0_in1[17]));
INVXL inst_cellmath__62_0_I308 (.Y(N830), .A(inst_cellmath__62_0_in1[18]));
INVXL inst_cellmath__62_0_I309 (.Y(N831), .A(inst_cellmath__62_0_in1[19]));
INVXL inst_cellmath__62_0_I310 (.Y(N832), .A(inst_cellmath__62_0_in1[20]));
INVXL inst_cellmath__62_0_I311 (.Y(N833), .A(inst_cellmath__62_0_in1[21]));
INVXL inst_cellmath__62_0_I312 (.Y(N834), .A(inst_cellmath__62_0_in1[22]));
INVXL inst_cellmath__62_0_I313 (.Y(N835), .A(inst_cellmath__62_0_in1[23]));
INVXL inst_cellmath__62_0_I314 (.Y(N836), .A(inst_cellmath__62_0_in1[24]));
INVXL inst_cellmath__62_0_I315 (.Y(N837), .A(inst_cellmath__62_0_in0[0]));
NOR2XL inst_cellmath__62_0_I49 (.Y(inst_cellmath__62_0_out1[4]), .A(N837), .B(N825));
NOR2XL inst_cellmath__62_0_I50 (.Y(inst_cellmath__62_0_out0[5]), .A(N837), .B(N826));
NOR2XL inst_cellmath__62_0_I51 (.Y(N313), .A(N837), .B(N827));
NOR2XL inst_cellmath__62_0_I52 (.Y(N315), .A(N837), .B(N828));
NOR2XL inst_cellmath__62_0_I53 (.Y(N317), .A(N837), .B(N829));
NOR2XL inst_cellmath__62_0_I54 (.Y(N319), .A(N837), .B(N830));
NOR2XL inst_cellmath__62_0_I55 (.Y(N321), .A(N837), .B(N831));
NOR2XL inst_cellmath__62_0_I56 (.Y(N323), .A(N837), .B(N832));
NOR2XL inst_cellmath__62_0_I57 (.Y(N325), .A(N837), .B(N833));
NOR2XL inst_cellmath__62_0_I58 (.Y(N327), .A(N837), .B(N834));
NOR2XL inst_cellmath__62_0_I59 (.Y(N329), .A(N837), .B(N835));
NOR2XL inst_cellmath__62_0_I60 (.Y(N331), .A(N837), .B(N836));
INVXL inst_cellmath__62_0_I316 (.Y(N838), .A(inst_cellmath__62_0_in0[1]));
NOR2XL inst_cellmath__62_0_I66 (.Y(inst_cellmath__62_0_out1[5]), .A(N838), .B(N825));
NOR2XL inst_cellmath__62_0_I67 (.Y(inst_cellmath__62_0_out1[6]), .A(N838), .B(N826));
NOR2XL inst_cellmath__62_0_I68 (.Y(N348), .A(N838), .B(N827));
NOR2XL inst_cellmath__62_0_I69 (.Y(N350), .A(N838), .B(N828));
NOR2XL inst_cellmath__62_0_I70 (.Y(N352), .A(N838), .B(N829));
NOR2XL inst_cellmath__62_0_I71 (.Y(N354), .A(N838), .B(N830));
NOR2XL inst_cellmath__62_0_I72 (.Y(N356), .A(N838), .B(N831));
NOR2XL inst_cellmath__62_0_I73 (.Y(N358), .A(N838), .B(N832));
NOR2XL inst_cellmath__62_0_I74 (.Y(N360), .A(N838), .B(N833));
NOR2XL inst_cellmath__62_0_I75 (.Y(N362), .A(N838), .B(N834));
NOR2XL inst_cellmath__62_0_I76 (.Y(N364), .A(N838), .B(N835));
NOR2XL inst_cellmath__62_0_I77 (.Y(N366), .A(N838), .B(N836));
INVXL inst_cellmath__62_0_I317 (.Y(N839), .A(inst_cellmath__62_0_in0[2]));
NOR2XL inst_cellmath__62_0_I83 (.Y(N379), .A(N839), .B(N825));
NOR2XL inst_cellmath__62_0_I84 (.Y(N381), .A(N839), .B(N826));
NOR2XL inst_cellmath__62_0_I85 (.Y(N383), .A(N839), .B(N827));
NOR2XL inst_cellmath__62_0_I86 (.Y(N385), .A(N839), .B(N828));
NOR2XL inst_cellmath__62_0_I87 (.Y(N387), .A(N839), .B(N829));
NOR2XL inst_cellmath__62_0_I88 (.Y(N389), .A(N839), .B(N830));
NOR2XL inst_cellmath__62_0_I89 (.Y(N391), .A(N839), .B(N831));
NOR2XL inst_cellmath__62_0_I90 (.Y(N393), .A(N839), .B(N832));
NOR2XL inst_cellmath__62_0_I91 (.Y(N395), .A(N839), .B(N833));
NOR2XL inst_cellmath__62_0_I92 (.Y(N397), .A(N839), .B(N834));
NOR2XL inst_cellmath__62_0_I93 (.Y(N399), .A(N839), .B(N835));
NOR2XL inst_cellmath__62_0_I94 (.Y(N401), .A(N839), .B(N836));
INVXL inst_cellmath__62_0_I318 (.Y(N840), .A(inst_cellmath__62_0_in0[3]));
NOR2XL inst_cellmath__62_0_I100 (.Y(N414), .A(N840), .B(N825));
NOR2XL inst_cellmath__62_0_I101 (.Y(N416), .A(N840), .B(N826));
NOR2XL inst_cellmath__62_0_I102 (.Y(N418), .A(N840), .B(N827));
NOR2XL inst_cellmath__62_0_I103 (.Y(N420), .A(N840), .B(N828));
NOR2XL inst_cellmath__62_0_I104 (.Y(N422), .A(N840), .B(N829));
NOR2XL inst_cellmath__62_0_I105 (.Y(N424), .A(N840), .B(N830));
NOR2XL inst_cellmath__62_0_I106 (.Y(N426), .A(N840), .B(N831));
NOR2XL inst_cellmath__62_0_I107 (.Y(N428), .A(N840), .B(N832));
NOR2XL inst_cellmath__62_0_I108 (.Y(N430), .A(N840), .B(N833));
NOR2XL inst_cellmath__62_0_I109 (.Y(N432), .A(N840), .B(N834));
NOR2XL inst_cellmath__62_0_I110 (.Y(N434), .A(N840), .B(N835));
NOR2XL inst_cellmath__62_0_I111 (.Y(N436), .A(N840), .B(N836));
INVXL inst_cellmath__62_0_I319 (.Y(N841), .A(inst_cellmath__62_0_in0[4]));
NOR2XL inst_cellmath__62_0_I117 (.Y(N449), .A(N841), .B(N825));
NOR2XL inst_cellmath__62_0_I118 (.Y(N451), .A(N841), .B(N826));
NOR2XL inst_cellmath__62_0_I119 (.Y(N453), .A(N841), .B(N827));
NOR2XL inst_cellmath__62_0_I120 (.Y(N455), .A(N841), .B(N828));
NOR2XL inst_cellmath__62_0_I121 (.Y(N457), .A(N841), .B(N829));
NOR2XL inst_cellmath__62_0_I122 (.Y(N459), .A(N841), .B(N830));
NOR2XL inst_cellmath__62_0_I123 (.Y(N461), .A(N841), .B(N831));
NOR2XL inst_cellmath__62_0_I124 (.Y(N463), .A(N841), .B(N832));
NOR2XL inst_cellmath__62_0_I125 (.Y(N465), .A(N841), .B(N833));
NOR2XL inst_cellmath__62_0_I126 (.Y(N467), .A(N841), .B(N834));
NOR2XL inst_cellmath__62_0_I127 (.Y(N469), .A(N841), .B(N835));
NOR2XL inst_cellmath__62_0_I128 (.Y(N471), .A(N841), .B(N836));
INVXL inst_cellmath__62_0_I320 (.Y(N842), .A(inst_cellmath__62_0_in0[5]));
NOR2XL inst_cellmath__62_0_I134 (.Y(N484), .A(N842), .B(N825));
NOR2XL inst_cellmath__62_0_I135 (.Y(N486), .A(N842), .B(N826));
NOR2XL inst_cellmath__62_0_I136 (.Y(N488), .A(N842), .B(N827));
NOR2XL inst_cellmath__62_0_I137 (.Y(N490), .A(N842), .B(N828));
NOR2XL inst_cellmath__62_0_I138 (.Y(N492), .A(N842), .B(N829));
NOR2XL inst_cellmath__62_0_I139 (.Y(N494), .A(N842), .B(N830));
NOR2XL inst_cellmath__62_0_I140 (.Y(N496), .A(N842), .B(N831));
NOR2XL inst_cellmath__62_0_I141 (.Y(N498), .A(N842), .B(N832));
NOR2XL inst_cellmath__62_0_I142 (.Y(N500), .A(N842), .B(N833));
NOR2XL inst_cellmath__62_0_I143 (.Y(N502), .A(N842), .B(N834));
NOR2XL inst_cellmath__62_0_I144 (.Y(N504), .A(N842), .B(N835));
NOR2XL inst_cellmath__62_0_I145 (.Y(N506), .A(N842), .B(N836));
INVXL inst_cellmath__62_0_I321 (.Y(N843), .A(inst_cellmath__62_0_in0[6]));
NOR2XL inst_cellmath__62_0_I151 (.Y(N519), .A(N843), .B(N825));
NOR2XL inst_cellmath__62_0_I152 (.Y(N521), .A(N843), .B(N826));
NOR2XL inst_cellmath__62_0_I153 (.Y(N523), .A(N843), .B(N827));
NOR2XL inst_cellmath__62_0_I154 (.Y(N525), .A(N843), .B(N828));
NOR2XL inst_cellmath__62_0_I155 (.Y(N527), .A(N843), .B(N829));
NOR2XL inst_cellmath__62_0_I156 (.Y(N529), .A(N843), .B(N830));
NOR2XL inst_cellmath__62_0_I157 (.Y(N531), .A(N843), .B(N831));
NOR2XL inst_cellmath__62_0_I158 (.Y(N533), .A(N843), .B(N832));
NOR2XL inst_cellmath__62_0_I159 (.Y(N535), .A(N843), .B(N833));
NOR2XL inst_cellmath__62_0_I160 (.Y(N537), .A(N843), .B(N834));
NOR2XL inst_cellmath__62_0_I161 (.Y(N539), .A(N843), .B(N835));
NOR2XL inst_cellmath__62_0_I162 (.Y(N541), .A(N843), .B(N836));
INVXL inst_cellmath__62_0_I322 (.Y(N844), .A(inst_cellmath__62_0_in0[7]));
NOR2XL inst_cellmath__62_0_I168 (.Y(N554), .A(N844), .B(N825));
NOR2XL inst_cellmath__62_0_I169 (.Y(N556), .A(N844), .B(N826));
NOR2XL inst_cellmath__62_0_I170 (.Y(N558), .A(N844), .B(N827));
NOR2XL inst_cellmath__62_0_I171 (.Y(N560), .A(N844), .B(N828));
NOR2XL inst_cellmath__62_0_I172 (.Y(N562), .A(N844), .B(N829));
NOR2XL inst_cellmath__62_0_I173 (.Y(N564), .A(N844), .B(N830));
NOR2XL inst_cellmath__62_0_I174 (.Y(N566), .A(N844), .B(N831));
NOR2XL inst_cellmath__62_0_I175 (.Y(N568), .A(N844), .B(N832));
NOR2XL inst_cellmath__62_0_I176 (.Y(N570), .A(N844), .B(N833));
NOR2XL inst_cellmath__62_0_I177 (.Y(N572), .A(N844), .B(N834));
NOR2XL inst_cellmath__62_0_I178 (.Y(N574), .A(N844), .B(N835));
NOR2XL inst_cellmath__62_0_I179 (.Y(N576), .A(N844), .B(N836));
INVXL inst_cellmath__62_0_I323 (.Y(N845), .A(inst_cellmath__62_0_in0[8]));
NOR2XL inst_cellmath__62_0_I185 (.Y(N589), .A(N845), .B(N825));
NOR2XL inst_cellmath__62_0_I186 (.Y(N591), .A(N845), .B(N826));
NOR2XL inst_cellmath__62_0_I187 (.Y(N593), .A(N845), .B(N827));
NOR2XL inst_cellmath__62_0_I188 (.Y(N595), .A(N845), .B(N828));
NOR2XL inst_cellmath__62_0_I189 (.Y(N597), .A(N845), .B(N829));
NOR2XL inst_cellmath__62_0_I190 (.Y(N599), .A(N845), .B(N830));
NOR2XL inst_cellmath__62_0_I191 (.Y(N601), .A(N845), .B(N831));
NOR2XL inst_cellmath__62_0_I192 (.Y(N603), .A(N845), .B(N832));
NOR2XL inst_cellmath__62_0_I193 (.Y(N605), .A(N845), .B(N833));
NOR2XL inst_cellmath__62_0_I194 (.Y(N607), .A(N845), .B(N834));
NOR2XL inst_cellmath__62_0_I195 (.Y(N609), .A(N845), .B(N835));
NOR2XL inst_cellmath__62_0_I196 (.Y(N611), .A(N845), .B(N836));
INVXL inst_cellmath__62_0_I324 (.Y(N846), .A(inst_cellmath__62_0_in0[9]));
NOR2XL inst_cellmath__62_0_I202 (.Y(N624), .A(N846), .B(N825));
NOR2XL inst_cellmath__62_0_I203 (.Y(N626), .A(N846), .B(N826));
NOR2XL inst_cellmath__62_0_I204 (.Y(N628), .A(N846), .B(N827));
NOR2XL inst_cellmath__62_0_I205 (.Y(N630), .A(N846), .B(N828));
NOR2XL inst_cellmath__62_0_I206 (.Y(N632), .A(N846), .B(N829));
NOR2XL inst_cellmath__62_0_I207 (.Y(N634), .A(N846), .B(N830));
NOR2XL inst_cellmath__62_0_I208 (.Y(N636), .A(N846), .B(N831));
NOR2XL inst_cellmath__62_0_I209 (.Y(N638), .A(N846), .B(N832));
NOR2XL inst_cellmath__62_0_I210 (.Y(N640), .A(N846), .B(N833));
NOR2XL inst_cellmath__62_0_I211 (.Y(N642), .A(N846), .B(N834));
NOR2XL inst_cellmath__62_0_I212 (.Y(N644), .A(N846), .B(N835));
NOR2XL inst_cellmath__62_0_I213 (.Y(inst_cellmath__62_0_out1[24]), .A(N846), .B(N836));
ADDHX1 inst_cellmath__62_0_I215 (.CO(N650), .S(inst_cellmath__62_0_out0[6]), .A(N379), .B(N313));
ADDHX1 inst_cellmath__62_0_I216 (.CO(N652), .S(inst_cellmath__62_0_out1[7]), .A(N414), .B(N315));
ADDFX1 inst_cellmath__62_0_I217 (.CO(N654), .S(inst_cellmath__62_0_out0[7]), .A(N348), .B(N381), .CI(N650));
ADDHX1 inst_cellmath__62_0_I218 (.CO(N656), .S(N655), .A(N449), .B(N350));
ADDFX1 inst_cellmath__62_0_I219 (.CO(N658), .S(inst_cellmath__62_0_out1[8]), .A(N317), .B(N416), .CI(N383));
ADDFX1 inst_cellmath__62_0_I220 (.CO(inst_cellmath__62_0_out1[9]), .S(inst_cellmath__62_0_out0[8]), .A(N655), .B(N652), .CI(N654));
ADDHX1 inst_cellmath__62_0_I221 (.CO(N662), .S(N661), .A(N484), .B(N385));
ADDFX1 inst_cellmath__62_0_I222 (.CO(N664), .S(N663), .A(N319), .B(N451), .CI(N418));
ADDFX1 inst_cellmath__62_0_I223 (.CO(N666), .S(N665), .A(N656), .B(N352), .CI(N661));
ADDFX1 inst_cellmath__62_0_I224 (.CO(inst_cellmath__62_0_out1[10]), .S(inst_cellmath__62_0_out0[9]), .A(N663), .B(N658), .CI(N665));
ADDHX1 inst_cellmath__62_0_I225 (.CO(N670), .S(N669), .A(N519), .B(N420));
ADDFX1 inst_cellmath__62_0_I226 (.CO(N672), .S(N671), .A(N354), .B(N486), .CI(N453));
ADDFX1 inst_cellmath__62_0_I227 (.CO(N674), .S(N673), .A(N321), .B(N387), .CI(N662));
ADDFX1 inst_cellmath__62_0_I228 (.CO(N676), .S(N675), .A(N664), .B(N669), .CI(N671));
ADDFX1 inst_cellmath__62_0_I229 (.CO(inst_cellmath__62_0_out1[11]), .S(inst_cellmath__62_0_out0[10]), .A(N673), .B(N666), .CI(N675));
ADDHX1 inst_cellmath__62_0_I230 (.CO(N680), .S(N679), .A(N554), .B(N455));
ADDFX1 inst_cellmath__62_0_I231 (.CO(N682), .S(N681), .A(N389), .B(N521), .CI(N488));
ADDFX1 inst_cellmath__62_0_I232 (.CO(N684), .S(N683), .A(N356), .B(N422), .CI(N323));
ADDFX1 inst_cellmath__62_0_I233 (.CO(N686), .S(N685), .A(N679), .B(N670), .CI(N672));
ADDFX1 inst_cellmath__62_0_I234 (.CO(N688), .S(N687), .A(N681), .B(N674), .CI(N683));
ADDFX1 inst_cellmath__62_0_I235 (.CO(inst_cellmath__62_0_out1[12]), .S(inst_cellmath__62_0_out0[11]), .A(N676), .B(N685), .CI(N687));
ADDHX1 inst_cellmath__62_0_I236 (.CO(N692), .S(N691), .A(N589), .B(N490));
ADDFX1 inst_cellmath__62_0_I237 (.CO(N694), .S(N693), .A(N424), .B(N556), .CI(N523));
ADDFX1 inst_cellmath__62_0_I238 (.CO(N696), .S(N695), .A(N391), .B(N457), .CI(N325));
ADDFX1 inst_cellmath__62_0_I239 (.CO(N698), .S(N697), .A(N680), .B(N358), .CI(N691));
ADDFX1 inst_cellmath__62_0_I240 (.CO(N700), .S(N699), .A(N684), .B(N682), .CI(N693));
ADDFX1 inst_cellmath__62_0_I241 (.CO(N702), .S(N701), .A(N695), .B(N686), .CI(N697));
ADDFX1 inst_cellmath__62_0_I242 (.CO(inst_cellmath__62_0_out1[13]), .S(inst_cellmath__62_0_out0[12]), .A(N699), .B(N688), .CI(N701));
ADDHX1 inst_cellmath__62_0_I243 (.CO(N706), .S(N705), .A(N624), .B(N525));
ADDFX1 inst_cellmath__62_0_I244 (.CO(N708), .S(N707), .A(N459), .B(N591), .CI(N558));
ADDFX1 inst_cellmath__62_0_I245 (.CO(N710), .S(N709), .A(N426), .B(N492), .CI(N360));
ADDFX1 inst_cellmath__62_0_I246 (.CO(N712), .S(N711), .A(N393), .B(N327), .CI(N692));
ADDFX1 inst_cellmath__62_0_I247 (.CO(N714), .S(N713), .A(N694), .B(N705), .CI(N696));
ADDFX1 inst_cellmath__62_0_I248 (.CO(N716), .S(N715), .A(N698), .B(N707), .CI(N709));
ADDFX1 inst_cellmath__62_0_I249 (.CO(N718), .S(N717), .A(N700), .B(N711), .CI(N713));
ADDFX1 inst_cellmath__62_0_I250 (.CO(inst_cellmath__62_0_out1[14]), .S(inst_cellmath__62_0_out0[13]), .A(N715), .B(N702), .CI(N717));
ADDFX1 inst_cellmath__62_0_I251 (.CO(N722), .S(N721), .A(N494), .B(N626), .CI(N593));
ADDFX1 inst_cellmath__62_0_I252 (.CO(N724), .S(N723), .A(N560), .B(N527), .CI(N461));
ADDFX1 inst_cellmath__62_0_I253 (.CO(N726), .S(N725), .A(N362), .B(N395), .CI(N428));
ADDFX1 inst_cellmath__62_0_I254 (.CO(N728), .S(N727), .A(N329), .B(N706), .CI(N708));
ADDFX1 inst_cellmath__62_0_I255 (.CO(N730), .S(N729), .A(N712), .B(N710), .CI(N721));
ADDFX1 inst_cellmath__62_0_I256 (.CO(N732), .S(N731), .A(N725), .B(N723), .CI(N714));
ADDFX1 inst_cellmath__62_0_I257 (.CO(N734), .S(N733), .A(N716), .B(N727), .CI(N729));
ADDFX1 inst_cellmath__62_0_I258 (.CO(inst_cellmath__62_0_out1[15]), .S(inst_cellmath__62_0_out0[14]), .A(N718), .B(N731), .CI(N733));
ADDFX1 inst_cellmath__62_0_I259 (.CO(N738), .S(N737), .A(N562), .B(N529), .CI(N595));
ADDFX1 inst_cellmath__62_0_I260 (.CO(N740), .S(N739), .A(N496), .B(N628), .CI(N430));
ADDFX1 inst_cellmath__62_0_I261 (.CO(N742), .S(N741), .A(N463), .B(N397), .CI(N364));
ADDFX1 inst_cellmath__62_0_I262 (.CO(N744), .S(N743), .A(N722), .B(N331), .CI(N724));
ADDFX1 inst_cellmath__62_0_I263 (.CO(N746), .S(N745), .A(N737), .B(N726), .CI(N728));
ADDFX1 inst_cellmath__62_0_I264 (.CO(N748), .S(N747), .A(N741), .B(N739), .CI(N730));
ADDFX1 inst_cellmath__62_0_I265 (.CO(N750), .S(N749), .A(N732), .B(N743), .CI(N745));
ADDFX1 inst_cellmath__62_0_I266 (.CO(inst_cellmath__62_0_out1[16]), .S(inst_cellmath__62_0_out0[15]), .A(N747), .B(N734), .CI(N749));
ADDHX1 inst_cellmath__62_0_I267 (.CO(N754), .S(N753), .A(N564), .B(N531));
ADDFX1 inst_cellmath__62_0_I268 (.CO(N756), .S(N755), .A(N630), .B(N597), .CI(N465));
ADDFX1 inst_cellmath__62_0_I269 (.CO(N758), .S(N757), .A(N498), .B(N432), .CI(N399));
ADDFX1 inst_cellmath__62_0_I270 (.CO(N760), .S(N759), .A(N753), .B(N366), .CI(N738));
ADDFX1 inst_cellmath__62_0_I271 (.CO(N762), .S(N761), .A(N742), .B(N740), .CI(N755));
ADDFX1 inst_cellmath__62_0_I272 (.CO(N764), .S(N763), .A(N757), .B(N744), .CI(N759));
ADDFX1 inst_cellmath__62_0_I273 (.CO(N766), .S(N765), .A(N761), .B(N746), .CI(N748));
ADDFX1 inst_cellmath__62_0_I274 (.CO(inst_cellmath__62_0_out1[17]), .S(inst_cellmath__62_0_out0[16]), .A(N750), .B(N763), .CI(N765));
ADDFX1 inst_cellmath__62_0_I275 (.CO(N770), .S(N769), .A(N632), .B(N599), .CI(N566));
ADDFX1 inst_cellmath__62_0_I276 (.CO(N772), .S(N771), .A(N467), .B(N500), .CI(N533));
ADDFX1 inst_cellmath__62_0_I277 (.CO(N774), .S(N773), .A(N401), .B(N434), .CI(N754));
ADDFX1 inst_cellmath__62_0_I278 (.CO(N776), .S(N775), .A(N758), .B(N756), .CI(N769));
ADDFX1 inst_cellmath__62_0_I279 (.CO(N778), .S(N777), .A(N771), .B(N760), .CI(N773));
ADDFX1 inst_cellmath__62_0_I280 (.CO(N780), .S(N779), .A(N775), .B(N762), .CI(N764));
ADDFX1 inst_cellmath__62_0_I281 (.CO(inst_cellmath__62_0_out1[18]), .S(inst_cellmath__62_0_out0[17]), .A(N766), .B(N777), .CI(N779));
ADDFX1 inst_cellmath__62_0_I282 (.CO(N784), .S(N783), .A(N601), .B(N634), .CI(N535));
ADDFX1 inst_cellmath__62_0_I283 (.CO(N786), .S(N785), .A(N568), .B(N502), .CI(N469));
ADDFX1 inst_cellmath__62_0_I284 (.CO(N788), .S(N787), .A(N770), .B(N436), .CI(N772));
ADDFX1 inst_cellmath__62_0_I285 (.CO(N790), .S(N789), .A(N783), .B(N774), .CI(N785));
ADDFX1 inst_cellmath__62_0_I286 (.CO(N792), .S(N791), .A(N787), .B(N776), .CI(N778));
ADDFX1 inst_cellmath__62_0_I287 (.CO(inst_cellmath__62_0_out1[19]), .S(inst_cellmath__62_0_out0[18]), .A(N780), .B(N789), .CI(N791));
ADDFX1 inst_cellmath__62_0_I288 (.CO(N796), .S(N795), .A(N570), .B(N636), .CI(N603));
ADDFX1 inst_cellmath__62_0_I289 (.CO(N798), .S(N797), .A(N504), .B(N537), .CI(N471));
ADDFX1 inst_cellmath__62_0_I290 (.CO(N800), .S(N799), .A(N786), .B(N784), .CI(N795));
ADDFX1 inst_cellmath__62_0_I291 (.CO(N802), .S(N801), .A(N788), .B(N797), .CI(N790));
ADDFX1 inst_cellmath__62_0_I292 (.CO(inst_cellmath__62_0_out1[20]), .S(inst_cellmath__62_0_out0[19]), .A(N792), .B(N799), .CI(N801));
ADDFX1 inst_cellmath__62_0_I293 (.CO(N806), .S(N805), .A(N572), .B(N605), .CI(N638));
ADDFX1 inst_cellmath__62_0_I294 (.CO(N808), .S(N807), .A(N506), .B(N539), .CI(N796));
ADDFX1 inst_cellmath__62_0_I295 (.CO(N810), .S(N809), .A(N805), .B(N798), .CI(N807));
ADDFX1 inst_cellmath__62_0_I296 (.CO(inst_cellmath__62_0_out1[21]), .S(inst_cellmath__62_0_out0[20]), .A(N802), .B(N800), .CI(N809));
ADDFX1 inst_cellmath__62_0_I297 (.CO(N814), .S(N813), .A(N607), .B(N640), .CI(N574));
ADDFX1 inst_cellmath__62_0_I298 (.CO(N816), .S(N815), .A(N806), .B(N541), .CI(N813));
ADDFX1 inst_cellmath__62_0_I299 (.CO(inst_cellmath__62_0_out0[22]), .S(inst_cellmath__62_0_out0[21]), .A(N815), .B(N808), .CI(N810));
ADDFX1 inst_cellmath__62_0_I300 (.CO(N820), .S(N819), .A(N609), .B(N642), .CI(N576));
ADDFX1 inst_cellmath__62_0_I301 (.CO(inst_cellmath__62_0_out0[23]), .S(inst_cellmath__62_0_out1[22]), .A(N819), .B(N814), .CI(N816));
ADDFX1 inst_cellmath__62_0_I302 (.CO(inst_cellmath__62_0_out0[24]), .S(inst_cellmath__62_0_out1[23]), .A(N611), .B(N644), .CI(N820));
assign inst_cellmath__62_0_out0[0] = 1'B0;
assign inst_cellmath__62_0_out0[1] = 1'B0;
assign inst_cellmath__62_0_out0[2] = 1'B0;
assign inst_cellmath__62_0_out0[3] = 1'B0;
assign inst_cellmath__62_0_out0[4] = 1'B0;
assign inst_cellmath__62_0_out0[25] = 1'B0;
assign inst_cellmath__62_0_out0[26] = 1'B0;
assign inst_cellmath__62_0_out0[27] = 1'B0;
assign inst_cellmath__62_0_out0[28] = 1'B0;
assign inst_cellmath__62_0_out0[29] = 1'B0;
assign inst_cellmath__62_0_out0[30] = 1'B0;
assign inst_cellmath__62_0_out0[31] = 1'B0;
assign inst_cellmath__62_0_out0[32] = 1'B0;
assign inst_cellmath__62_0_out0[33] = 1'B0;
assign inst_cellmath__62_0_out0[34] = 1'B0;
assign inst_cellmath__62_0_out0[35] = 1'B0;
assign inst_cellmath__62_0_out0[36] = 1'B0;
assign inst_cellmath__62_0_out0[37] = 1'B0;
assign inst_cellmath__62_0_out0[38] = 1'B0;
assign inst_cellmath__62_0_out0[39] = 1'B0;
assign inst_cellmath__62_0_out1[0] = 1'B0;
assign inst_cellmath__62_0_out1[1] = 1'B0;
assign inst_cellmath__62_0_out1[2] = 1'B0;
assign inst_cellmath__62_0_out1[3] = 1'B0;
assign inst_cellmath__62_0_out1[25] = 1'B0;
assign inst_cellmath__62_0_out1[26] = 1'B0;
assign inst_cellmath__62_0_out1[27] = 1'B0;
assign inst_cellmath__62_0_out1[28] = 1'B0;
assign inst_cellmath__62_0_out1[29] = 1'B0;
assign inst_cellmath__62_0_out1[30] = 1'B0;
assign inst_cellmath__62_0_out1[31] = 1'B0;
assign inst_cellmath__62_0_out1[32] = 1'B0;
assign inst_cellmath__62_0_out1[33] = 1'B0;
assign inst_cellmath__62_0_out1[34] = 1'B0;
assign inst_cellmath__62_0_out1[35] = 1'B0;
assign inst_cellmath__62_0_out1[36] = 1'B0;
assign inst_cellmath__62_0_out1[37] = 1'B0;
assign inst_cellmath__62_0_out1[38] = 1'B0;
assign inst_cellmath__62_0_out1[39] = 1'B0;
endmodule

module cynw_cm_float_rcp_inst_cellmath__63_0_bdw1412651405_bdw (
	inst_cellmath__63_0_out0,
	inst_cellmath__63_0_out1,
	inst_cellmath__63_0_in0,
	inst_cellmath__63_0_in1,
	inst_cellmath__63_0_in2
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__63_0_out0,
	inst_cellmath__63_0_out1;
input [27:10] inst_cellmath__63_0_in0;
input  inst_cellmath__63_0_in1;
input [14:0] inst_cellmath__63_0_in2;
wire N414,N416,N418,N420,N422,N424,N426 
	,N428,N430,N432,N434,N436,N438,N440,N442 
	,N444,N462,N464,N466,N468,N470,N472,N474 
	,N476,N478,N480,N482,N484,N486,N488,N490 
	,N492,N506,N508,N510,N512,N514,N516,N518 
	,N520,N522,N524,N526,N528,N530,N532,N534 
	,N536,N538,N540,N554,N556,N558,N560,N562 
	,N564,N566,N568,N570,N572,N574,N576,N578 
	,N580,N582,N584,N586,N588,N602,N604,N606 
	,N608,N610,N612,N614,N616,N618,N620,N622 
	,N624,N626,N628,N630,N632,N634,N636,N650 
	,N652,N654,N656,N658,N660,N662,N664,N666 
	,N668,N670,N672,N674,N676,N678,N680,N682 
	,N684,N698,N700,N702,N704,N706,N708,N710 
	,N712,N714,N716,N718,N720,N722,N724,N726 
	,N728,N730,N732,N746,N748,N750,N752,N754 
	,N756,N758,N760,N762,N764,N766,N768,N770 
	,N772,N774,N776,N778,N780,N794,N796,N798 
	,N800,N802,N804,N806,N808,N810,N812,N814 
	,N816,N818,N820,N822,N824,N826,N828,N842 
	,N844,N846,N848,N850,N852,N854,N856,N858 
	,N860,N862,N864,N866,N868,N870,N872,N874 
	,N876,N890,N892,N894,N896,N898,N900,N902 
	,N904,N906,N908,N910,N912,N914,N916,N918 
	,N920,N922,N924,N938,N940,N942,N944,N946 
	,N948,N950,N952,N954,N956,N958,N960,N962 
	,N964,N966,N968,N970,N972,N986,N988,N990 
	,N992,N994,N996,N998,N1000,N1002,N1004,N1006 
	,N1008,N1010,N1012,N1014,N1016,N1018,N1020,N1034 
	,N1036,N1038,N1040,N1042,N1044,N1046,N1048,N1050 
	,N1052,N1054,N1056,N1058,N1060,N1062,N1064,N1066 
	,N1068,N1082,N1084,N1086,N1088,N1090,N1092,N1094 
	,N1096,N1098,N1100,N1102,N1104,N1106,N1108,N1110 
	,N1112,N1114,N1116,N1130,N1132,N1134,N1136,N1138 
	,N1140,N1142,N1144,N1146,N1148,N1150,N1152,N1154 
	,N1156,N1158,N1160,N1162,N1164,N1185,N1187,N1189 
	,N1190,N1191,N1193,N1196,N1197,N1198,N1199,N1200 
	,N1201,N1204,N1205,N1206,N1207,N1208,N1209,N1210 
	,N1211,N1214,N1215,N1216,N1217,N1218,N1219,N1220 
	,N1221,N1222,N1223,N1226,N1227,N1228,N1229,N1230 
	,N1231,N1232,N1233,N1234,N1235,N1236,N1237,N1240 
	,N1241,N1242,N1243,N1244,N1245,N1246,N1247,N1248 
	,N1249,N1250,N1251,N1252,N1253,N1256,N1257,N1258 
	,N1259,N1260,N1261,N1262,N1263,N1264,N1265,N1266 
	,N1267,N1268,N1269,N1270,N1271,N1274,N1275,N1276 
	,N1277,N1278,N1279,N1280,N1281,N1282,N1283,N1284 
	,N1285,N1286,N1287,N1288,N1289,N1290,N1291,N1294 
	,N1295,N1296,N1297,N1298,N1299,N1300,N1301,N1302 
	,N1303,N1304,N1305,N1306,N1307,N1308,N1309,N1310 
	,N1311,N1312,N1313,N1316,N1317,N1318,N1319,N1320 
	,N1321,N1322,N1323,N1324,N1325,N1326,N1327,N1328 
	,N1329,N1330,N1331,N1332,N1333,N1334,N1335,N1336 
	,N1337,N1340,N1341,N1342,N1343,N1344,N1345,N1346 
	,N1347,N1348,N1349,N1350,N1351,N1352,N1353,N1354 
	,N1355,N1356,N1357,N1358,N1359,N1360,N1361,N1362 
	,N1363,N1366,N1367,N1370,N1371,N1372,N1373,N1374 
	,N1375,N1376,N1377,N1378,N1379,N1380,N1381,N1382 
	,N1383,N1384,N1385,N1386,N1387,N1388,N1389,N1390 
	,N1391,N1392,N1393,N1396,N1397,N1398,N1399,N1400 
	,N1401,N1402,N1403,N1404,N1405,N1406,N1407,N1408 
	,N1409,N1410,N1411,N1412,N1413,N1414,N1415,N1416 
	,N1417,N1418,N1419,N1420,N1421,N1424,N1425,N1426 
	,N1427,N1428,N1429,N1430,N1431,N1432,N1433,N1434 
	,N1435,N1436,N1437,N1438,N1439,N1440,N1441,N1442 
	,N1443,N1444,N1445,N1446,N1447,N1448,N1449,N1452 
	,N1453,N1456,N1457,N1458,N1459,N1460,N1461,N1462 
	,N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470 
	,N1471,N1472,N1473,N1474,N1475,N1476,N1477,N1478 
	,N1479,N1482,N1483,N1484,N1485,N1486,N1487,N1488 
	,N1489,N1490,N1491,N1492,N1493,N1494,N1495,N1496 
	,N1497,N1498,N1499,N1500,N1501,N1502,N1503,N1504 
	,N1505,N1506,N1507,N1510,N1511,N1512,N1513,N1514 
	,N1515,N1516,N1517,N1518,N1519,N1520,N1521,N1522 
	,N1523,N1524,N1525,N1526,N1527,N1528,N1529,N1530 
	,N1531,N1532,N1533,N1536,N1537,N1538,N1539,N1540 
	,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548 
	,N1549,N1550,N1551,N1552,N1553,N1554,N1555,N1556 
	,N1557,N1560,N1561,N1562,N1563,N1564,N1565,N1566 
	,N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574 
	,N1575,N1576,N1577,N1578,N1579,N1582,N1583,N1584 
	,N1585,N1586,N1587,N1588,N1589,N1590,N1591,N1592 
	,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1602 
	,N1603,N1604,N1605,N1606,N1607,N1608,N1609,N1610 
	,N1611,N1612,N1613,N1614,N1615,N1616,N1617,N1620 
	,N1621,N1622,N1623,N1624,N1625,N1626,N1627,N1628 
	,N1629,N1630,N1631,N1632,N1633,N1636,N1637,N1638 
	,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646 
	,N1647,N1650,N1651,N1652,N1653,N1654,N1655,N1656 
	,N1657,N1658,N1659,N1662,N1663,N1664,N1665,N1666 
	,N1667,N1668,N1669,N1672,N1673,N1674,N1675,N1676 
	,N1677,N1680,N1681,N1682,N1683,N1686,N1687,N1803 
	,N1813,N1820,N1827,N1834,N1841,N1848,N1855,N1862 
	,N1869,N1876,N1883,N1890,N1897,N1904,N1911,N1918 
	,N1925,N1932,N1938,N1944,N1950,N1956,N1962,N1968 
	,N1974,N1980,N1986,N1992,N1998,N2004,N2010,N2016 
	,N2022;
INVXL inst_cellmath__63_0_I726 (.Y(N1813), .A(inst_cellmath__63_0_in0[10]));
INVXL inst_cellmath__63_0_I733 (.Y(N1820), .A(inst_cellmath__63_0_in0[11]));
INVXL inst_cellmath__63_0_I740 (.Y(N1827), .A(inst_cellmath__63_0_in0[12]));
INVXL inst_cellmath__63_0_I747 (.Y(N1834), .A(inst_cellmath__63_0_in0[13]));
INVXL inst_cellmath__63_0_I754 (.Y(N1841), .A(inst_cellmath__63_0_in0[14]));
INVXL inst_cellmath__63_0_I761 (.Y(N1848), .A(inst_cellmath__63_0_in0[15]));
INVXL inst_cellmath__63_0_I768 (.Y(N1855), .A(inst_cellmath__63_0_in0[16]));
INVXL inst_cellmath__63_0_I775 (.Y(N1862), .A(inst_cellmath__63_0_in0[17]));
INVXL inst_cellmath__63_0_I782 (.Y(N1869), .A(inst_cellmath__63_0_in0[18]));
INVXL inst_cellmath__63_0_I789 (.Y(N1876), .A(inst_cellmath__63_0_in0[19]));
INVXL inst_cellmath__63_0_I796 (.Y(N1883), .A(inst_cellmath__63_0_in0[20]));
INVXL inst_cellmath__63_0_I803 (.Y(N1890), .A(inst_cellmath__63_0_in0[21]));
INVXL inst_cellmath__63_0_I810 (.Y(N1897), .A(inst_cellmath__63_0_in0[22]));
INVXL inst_cellmath__63_0_I817 (.Y(N1904), .A(inst_cellmath__63_0_in0[23]));
INVXL inst_cellmath__63_0_I824 (.Y(N1911), .A(inst_cellmath__63_0_in0[24]));
INVXL inst_cellmath__63_0_I831 (.Y(N1918), .A(inst_cellmath__63_0_in0[25]));
INVXL inst_cellmath__63_0_I838 (.Y(N1925), .A(inst_cellmath__63_0_in0[26]));
INVXL inst_cellmath__63_0_I845 (.Y(N1932), .A(inst_cellmath__63_0_in0[27]));
INVXL inst_cellmath__63_0_I1002 (.Y(N1938), .A(inst_cellmath__63_0_in2[0]));
NOR2XL inst_cellmath__63_0_I66 (.Y(inst_cellmath__63_0_out1[0]), .A(N1938), .B(N1813));
NOR2XL inst_cellmath__63_0_I67 (.Y(inst_cellmath__63_0_out0[1]), .A(N1938), .B(N1820));
NOR2XL inst_cellmath__63_0_I68 (.Y(N414), .A(N1938), .B(N1827));
NOR2XL inst_cellmath__63_0_I69 (.Y(N416), .A(N1938), .B(N1834));
NOR2XL inst_cellmath__63_0_I70 (.Y(N418), .A(N1938), .B(N1841));
NOR2XL inst_cellmath__63_0_I71 (.Y(N420), .A(N1938), .B(N1848));
NOR2XL inst_cellmath__63_0_I72 (.Y(N422), .A(N1938), .B(N1855));
NOR2XL inst_cellmath__63_0_I73 (.Y(N424), .A(N1938), .B(N1862));
NOR2XL inst_cellmath__63_0_I74 (.Y(N426), .A(N1938), .B(N1869));
NOR2XL inst_cellmath__63_0_I75 (.Y(N428), .A(N1938), .B(N1876));
NOR2XL inst_cellmath__63_0_I76 (.Y(N430), .A(N1938), .B(N1883));
NOR2XL inst_cellmath__63_0_I77 (.Y(N432), .A(N1938), .B(N1890));
NOR2XL inst_cellmath__63_0_I78 (.Y(N434), .A(N1938), .B(N1897));
NOR2XL inst_cellmath__63_0_I79 (.Y(N436), .A(N1938), .B(N1904));
NOR2XL inst_cellmath__63_0_I80 (.Y(N438), .A(N1938), .B(N1911));
NOR2XL inst_cellmath__63_0_I81 (.Y(N440), .A(N1938), .B(N1918));
NOR2XL inst_cellmath__63_0_I82 (.Y(N442), .A(N1938), .B(N1925));
NOR2XL inst_cellmath__63_0_I83 (.Y(N444), .A(N1938), .B(N1932));
INVXL inst_cellmath__63_0_I1003 (.Y(N1944), .A(inst_cellmath__63_0_in2[1]));
NOR2XL inst_cellmath__63_0_I89 (.Y(inst_cellmath__63_0_out1[1]), .A(N1944), .B(N1813));
NOR2XL inst_cellmath__63_0_I90 (.Y(inst_cellmath__63_0_out1[2]), .A(N1944), .B(N1820));
NOR2XL inst_cellmath__63_0_I91 (.Y(N462), .A(N1944), .B(N1827));
NOR2XL inst_cellmath__63_0_I92 (.Y(N464), .A(N1944), .B(N1834));
NOR2XL inst_cellmath__63_0_I93 (.Y(N466), .A(N1944), .B(N1841));
NOR2XL inst_cellmath__63_0_I94 (.Y(N468), .A(N1944), .B(N1848));
NOR2XL inst_cellmath__63_0_I95 (.Y(N470), .A(N1944), .B(N1855));
NOR2XL inst_cellmath__63_0_I96 (.Y(N472), .A(N1944), .B(N1862));
NOR2XL inst_cellmath__63_0_I97 (.Y(N474), .A(N1944), .B(N1869));
NOR2XL inst_cellmath__63_0_I98 (.Y(N476), .A(N1944), .B(N1876));
NOR2XL inst_cellmath__63_0_I99 (.Y(N478), .A(N1944), .B(N1883));
NOR2XL inst_cellmath__63_0_I100 (.Y(N480), .A(N1944), .B(N1890));
NOR2XL inst_cellmath__63_0_I101 (.Y(N482), .A(N1944), .B(N1897));
NOR2XL inst_cellmath__63_0_I102 (.Y(N484), .A(N1944), .B(N1904));
NOR2XL inst_cellmath__63_0_I103 (.Y(N486), .A(N1944), .B(N1911));
NOR2XL inst_cellmath__63_0_I104 (.Y(N488), .A(N1944), .B(N1918));
NOR2XL inst_cellmath__63_0_I105 (.Y(N490), .A(N1944), .B(N1925));
NOR2XL inst_cellmath__63_0_I106 (.Y(N492), .A(N1944), .B(N1932));
INVXL inst_cellmath__63_0_I1004 (.Y(N1950), .A(inst_cellmath__63_0_in2[2]));
NOR2XL inst_cellmath__63_0_I112 (.Y(N506), .A(N1950), .B(N1813));
NOR2XL inst_cellmath__63_0_I113 (.Y(N508), .A(N1950), .B(N1820));
NOR2XL inst_cellmath__63_0_I114 (.Y(N510), .A(N1950), .B(N1827));
NOR2XL inst_cellmath__63_0_I115 (.Y(N512), .A(N1950), .B(N1834));
NOR2XL inst_cellmath__63_0_I116 (.Y(N514), .A(N1950), .B(N1841));
NOR2XL inst_cellmath__63_0_I117 (.Y(N516), .A(N1950), .B(N1848));
NOR2XL inst_cellmath__63_0_I118 (.Y(N518), .A(N1950), .B(N1855));
NOR2XL inst_cellmath__63_0_I119 (.Y(N520), .A(N1950), .B(N1862));
NOR2XL inst_cellmath__63_0_I120 (.Y(N522), .A(N1950), .B(N1869));
NOR2XL inst_cellmath__63_0_I121 (.Y(N524), .A(N1950), .B(N1876));
NOR2XL inst_cellmath__63_0_I122 (.Y(N526), .A(N1950), .B(N1883));
NOR2XL inst_cellmath__63_0_I123 (.Y(N528), .A(N1950), .B(N1890));
NOR2XL inst_cellmath__63_0_I124 (.Y(N530), .A(N1950), .B(N1897));
NOR2XL inst_cellmath__63_0_I125 (.Y(N532), .A(N1950), .B(N1904));
NOR2XL inst_cellmath__63_0_I126 (.Y(N534), .A(N1950), .B(N1911));
NOR2XL inst_cellmath__63_0_I127 (.Y(N536), .A(N1950), .B(N1918));
NOR2XL inst_cellmath__63_0_I128 (.Y(N538), .A(N1950), .B(N1925));
NOR2XL inst_cellmath__63_0_I129 (.Y(N540), .A(N1950), .B(N1932));
INVXL inst_cellmath__63_0_I1005 (.Y(N1956), .A(inst_cellmath__63_0_in2[3]));
NOR2XL inst_cellmath__63_0_I135 (.Y(N554), .A(N1956), .B(N1813));
NOR2XL inst_cellmath__63_0_I136 (.Y(N556), .A(N1956), .B(N1820));
NOR2XL inst_cellmath__63_0_I137 (.Y(N558), .A(N1956), .B(N1827));
NOR2XL inst_cellmath__63_0_I138 (.Y(N560), .A(N1956), .B(N1834));
NOR2XL inst_cellmath__63_0_I139 (.Y(N562), .A(N1956), .B(N1841));
NOR2XL inst_cellmath__63_0_I140 (.Y(N564), .A(N1956), .B(N1848));
NOR2XL inst_cellmath__63_0_I141 (.Y(N566), .A(N1956), .B(N1855));
NOR2XL inst_cellmath__63_0_I142 (.Y(N568), .A(N1956), .B(N1862));
NOR2XL inst_cellmath__63_0_I143 (.Y(N570), .A(N1956), .B(N1869));
NOR2XL inst_cellmath__63_0_I144 (.Y(N572), .A(N1956), .B(N1876));
NOR2XL inst_cellmath__63_0_I145 (.Y(N574), .A(N1956), .B(N1883));
NOR2XL inst_cellmath__63_0_I146 (.Y(N576), .A(N1956), .B(N1890));
NOR2XL inst_cellmath__63_0_I147 (.Y(N578), .A(N1956), .B(N1897));
NOR2XL inst_cellmath__63_0_I148 (.Y(N580), .A(N1956), .B(N1904));
NOR2XL inst_cellmath__63_0_I149 (.Y(N582), .A(N1956), .B(N1911));
NOR2XL inst_cellmath__63_0_I150 (.Y(N584), .A(N1956), .B(N1918));
NOR2XL inst_cellmath__63_0_I151 (.Y(N586), .A(N1956), .B(N1925));
NOR2XL inst_cellmath__63_0_I152 (.Y(N588), .A(N1956), .B(N1932));
INVXL inst_cellmath__63_0_I1006 (.Y(N1962), .A(inst_cellmath__63_0_in2[4]));
NOR2XL inst_cellmath__63_0_I158 (.Y(N602), .A(N1962), .B(N1813));
NOR2XL inst_cellmath__63_0_I159 (.Y(N604), .A(N1962), .B(N1820));
NOR2XL inst_cellmath__63_0_I160 (.Y(N606), .A(N1962), .B(N1827));
NOR2XL inst_cellmath__63_0_I161 (.Y(N608), .A(N1962), .B(N1834));
NOR2XL inst_cellmath__63_0_I162 (.Y(N610), .A(N1962), .B(N1841));
NOR2XL inst_cellmath__63_0_I163 (.Y(N612), .A(N1962), .B(N1848));
NOR2XL inst_cellmath__63_0_I164 (.Y(N614), .A(N1962), .B(N1855));
NOR2XL inst_cellmath__63_0_I165 (.Y(N616), .A(N1962), .B(N1862));
NOR2XL inst_cellmath__63_0_I166 (.Y(N618), .A(N1962), .B(N1869));
NOR2XL inst_cellmath__63_0_I167 (.Y(N620), .A(N1962), .B(N1876));
NOR2XL inst_cellmath__63_0_I168 (.Y(N622), .A(N1962), .B(N1883));
NOR2XL inst_cellmath__63_0_I169 (.Y(N624), .A(N1962), .B(N1890));
NOR2XL inst_cellmath__63_0_I170 (.Y(N626), .A(N1962), .B(N1897));
NOR2XL inst_cellmath__63_0_I171 (.Y(N628), .A(N1962), .B(N1904));
NOR2XL inst_cellmath__63_0_I172 (.Y(N630), .A(N1962), .B(N1911));
NOR2XL inst_cellmath__63_0_I173 (.Y(N632), .A(N1962), .B(N1918));
NOR2XL inst_cellmath__63_0_I174 (.Y(N634), .A(N1962), .B(N1925));
NOR2XL inst_cellmath__63_0_I175 (.Y(N636), .A(N1962), .B(N1932));
INVXL inst_cellmath__63_0_I1007 (.Y(N1968), .A(inst_cellmath__63_0_in2[5]));
NOR2XL inst_cellmath__63_0_I181 (.Y(N650), .A(N1968), .B(N1813));
NOR2XL inst_cellmath__63_0_I182 (.Y(N652), .A(N1968), .B(N1820));
NOR2XL inst_cellmath__63_0_I183 (.Y(N654), .A(N1968), .B(N1827));
NOR2XL inst_cellmath__63_0_I184 (.Y(N656), .A(N1968), .B(N1834));
NOR2XL inst_cellmath__63_0_I185 (.Y(N658), .A(N1968), .B(N1841));
NOR2XL inst_cellmath__63_0_I186 (.Y(N660), .A(N1968), .B(N1848));
NOR2XL inst_cellmath__63_0_I187 (.Y(N662), .A(N1968), .B(N1855));
NOR2XL inst_cellmath__63_0_I188 (.Y(N664), .A(N1968), .B(N1862));
NOR2XL inst_cellmath__63_0_I189 (.Y(N666), .A(N1968), .B(N1869));
NOR2XL inst_cellmath__63_0_I190 (.Y(N668), .A(N1968), .B(N1876));
NOR2XL inst_cellmath__63_0_I191 (.Y(N670), .A(N1968), .B(N1883));
NOR2XL inst_cellmath__63_0_I192 (.Y(N672), .A(N1968), .B(N1890));
NOR2XL inst_cellmath__63_0_I193 (.Y(N674), .A(N1968), .B(N1897));
NOR2XL inst_cellmath__63_0_I194 (.Y(N676), .A(N1968), .B(N1904));
NOR2XL inst_cellmath__63_0_I195 (.Y(N678), .A(N1968), .B(N1911));
NOR2XL inst_cellmath__63_0_I196 (.Y(N680), .A(N1968), .B(N1918));
NOR2XL inst_cellmath__63_0_I197 (.Y(N682), .A(N1968), .B(N1925));
NOR2XL inst_cellmath__63_0_I198 (.Y(N684), .A(N1968), .B(N1932));
INVXL inst_cellmath__63_0_I1008 (.Y(N1974), .A(inst_cellmath__63_0_in2[6]));
NOR2XL inst_cellmath__63_0_I204 (.Y(N698), .A(N1974), .B(N1813));
NOR2XL inst_cellmath__63_0_I205 (.Y(N700), .A(N1974), .B(N1820));
NOR2XL inst_cellmath__63_0_I206 (.Y(N702), .A(N1974), .B(N1827));
NOR2XL inst_cellmath__63_0_I207 (.Y(N704), .A(N1974), .B(N1834));
NOR2XL inst_cellmath__63_0_I208 (.Y(N706), .A(N1974), .B(N1841));
NOR2XL inst_cellmath__63_0_I209 (.Y(N708), .A(N1974), .B(N1848));
NOR2XL inst_cellmath__63_0_I210 (.Y(N710), .A(N1974), .B(N1855));
NOR2XL inst_cellmath__63_0_I211 (.Y(N712), .A(N1974), .B(N1862));
NOR2XL inst_cellmath__63_0_I212 (.Y(N714), .A(N1974), .B(N1869));
NOR2XL inst_cellmath__63_0_I213 (.Y(N716), .A(N1974), .B(N1876));
NOR2XL inst_cellmath__63_0_I214 (.Y(N718), .A(N1974), .B(N1883));
NOR2XL inst_cellmath__63_0_I215 (.Y(N720), .A(N1974), .B(N1890));
NOR2XL inst_cellmath__63_0_I216 (.Y(N722), .A(N1974), .B(N1897));
NOR2XL inst_cellmath__63_0_I217 (.Y(N724), .A(N1974), .B(N1904));
NOR2XL inst_cellmath__63_0_I218 (.Y(N726), .A(N1974), .B(N1911));
NOR2XL inst_cellmath__63_0_I219 (.Y(N728), .A(N1974), .B(N1918));
NOR2XL inst_cellmath__63_0_I220 (.Y(N730), .A(N1974), .B(N1925));
NOR2XL inst_cellmath__63_0_I221 (.Y(N732), .A(N1974), .B(N1932));
INVXL inst_cellmath__63_0_I1009 (.Y(N1980), .A(inst_cellmath__63_0_in2[7]));
NOR2XL inst_cellmath__63_0_I227 (.Y(N746), .A(N1980), .B(N1813));
NOR2XL inst_cellmath__63_0_I228 (.Y(N748), .A(N1980), .B(N1820));
NOR2XL inst_cellmath__63_0_I229 (.Y(N750), .A(N1980), .B(N1827));
NOR2XL inst_cellmath__63_0_I230 (.Y(N752), .A(N1980), .B(N1834));
NOR2XL inst_cellmath__63_0_I231 (.Y(N754), .A(N1980), .B(N1841));
NOR2XL inst_cellmath__63_0_I232 (.Y(N756), .A(N1980), .B(N1848));
NOR2XL inst_cellmath__63_0_I233 (.Y(N758), .A(N1980), .B(N1855));
NOR2XL inst_cellmath__63_0_I234 (.Y(N760), .A(N1980), .B(N1862));
NOR2XL inst_cellmath__63_0_I235 (.Y(N762), .A(N1980), .B(N1869));
NOR2XL inst_cellmath__63_0_I236 (.Y(N764), .A(N1980), .B(N1876));
NOR2XL inst_cellmath__63_0_I237 (.Y(N766), .A(N1980), .B(N1883));
NOR2XL inst_cellmath__63_0_I238 (.Y(N768), .A(N1980), .B(N1890));
NOR2XL inst_cellmath__63_0_I239 (.Y(N770), .A(N1980), .B(N1897));
NOR2XL inst_cellmath__63_0_I240 (.Y(N772), .A(N1980), .B(N1904));
NOR2XL inst_cellmath__63_0_I241 (.Y(N774), .A(N1980), .B(N1911));
NOR2XL inst_cellmath__63_0_I242 (.Y(N776), .A(N1980), .B(N1918));
NOR2XL inst_cellmath__63_0_I243 (.Y(N778), .A(N1980), .B(N1925));
NOR2XL inst_cellmath__63_0_I244 (.Y(N780), .A(N1980), .B(N1932));
INVXL inst_cellmath__63_0_I1010 (.Y(N1986), .A(inst_cellmath__63_0_in2[8]));
NOR2XL inst_cellmath__63_0_I250 (.Y(N794), .A(N1986), .B(N1813));
NOR2XL inst_cellmath__63_0_I251 (.Y(N796), .A(N1986), .B(N1820));
NOR2XL inst_cellmath__63_0_I252 (.Y(N798), .A(N1986), .B(N1827));
NOR2XL inst_cellmath__63_0_I253 (.Y(N800), .A(N1986), .B(N1834));
NOR2XL inst_cellmath__63_0_I254 (.Y(N802), .A(N1986), .B(N1841));
NOR2XL inst_cellmath__63_0_I255 (.Y(N804), .A(N1986), .B(N1848));
NOR2XL inst_cellmath__63_0_I256 (.Y(N806), .A(N1986), .B(N1855));
NOR2XL inst_cellmath__63_0_I257 (.Y(N808), .A(N1986), .B(N1862));
NOR2XL inst_cellmath__63_0_I258 (.Y(N810), .A(N1986), .B(N1869));
NOR2XL inst_cellmath__63_0_I259 (.Y(N812), .A(N1986), .B(N1876));
NOR2XL inst_cellmath__63_0_I260 (.Y(N814), .A(N1986), .B(N1883));
NOR2XL inst_cellmath__63_0_I261 (.Y(N816), .A(N1986), .B(N1890));
NOR2XL inst_cellmath__63_0_I262 (.Y(N818), .A(N1986), .B(N1897));
NOR2XL inst_cellmath__63_0_I263 (.Y(N820), .A(N1986), .B(N1904));
NOR2XL inst_cellmath__63_0_I264 (.Y(N822), .A(N1986), .B(N1911));
NOR2XL inst_cellmath__63_0_I265 (.Y(N824), .A(N1986), .B(N1918));
NOR2XL inst_cellmath__63_0_I266 (.Y(N826), .A(N1986), .B(N1925));
NOR2XL inst_cellmath__63_0_I267 (.Y(N828), .A(N1986), .B(N1932));
INVXL inst_cellmath__63_0_I1011 (.Y(N1992), .A(inst_cellmath__63_0_in2[9]));
NOR2XL inst_cellmath__63_0_I273 (.Y(N842), .A(N1992), .B(N1813));
NOR2XL inst_cellmath__63_0_I274 (.Y(N844), .A(N1992), .B(N1820));
NOR2XL inst_cellmath__63_0_I275 (.Y(N846), .A(N1992), .B(N1827));
NOR2XL inst_cellmath__63_0_I276 (.Y(N848), .A(N1992), .B(N1834));
NOR2XL inst_cellmath__63_0_I277 (.Y(N850), .A(N1992), .B(N1841));
NOR2XL inst_cellmath__63_0_I278 (.Y(N852), .A(N1992), .B(N1848));
NOR2XL inst_cellmath__63_0_I279 (.Y(N854), .A(N1992), .B(N1855));
NOR2XL inst_cellmath__63_0_I280 (.Y(N856), .A(N1992), .B(N1862));
NOR2XL inst_cellmath__63_0_I281 (.Y(N858), .A(N1992), .B(N1869));
NOR2XL inst_cellmath__63_0_I282 (.Y(N860), .A(N1992), .B(N1876));
NOR2XL inst_cellmath__63_0_I283 (.Y(N862), .A(N1992), .B(N1883));
NOR2XL inst_cellmath__63_0_I284 (.Y(N864), .A(N1992), .B(N1890));
NOR2XL inst_cellmath__63_0_I285 (.Y(N866), .A(N1992), .B(N1897));
NOR2XL inst_cellmath__63_0_I286 (.Y(N868), .A(N1992), .B(N1904));
NOR2XL inst_cellmath__63_0_I287 (.Y(N870), .A(N1992), .B(N1911));
NOR2XL inst_cellmath__63_0_I288 (.Y(N872), .A(N1992), .B(N1918));
NOR2XL inst_cellmath__63_0_I289 (.Y(N874), .A(N1992), .B(N1925));
NOR2XL inst_cellmath__63_0_I290 (.Y(N876), .A(N1992), .B(N1932));
INVXL inst_cellmath__63_0_I1012 (.Y(N1998), .A(inst_cellmath__63_0_in2[10]));
NOR2XL inst_cellmath__63_0_I296 (.Y(N890), .A(N1998), .B(N1813));
NOR2XL inst_cellmath__63_0_I297 (.Y(N892), .A(N1998), .B(N1820));
NOR2XL inst_cellmath__63_0_I298 (.Y(N894), .A(N1998), .B(N1827));
NOR2XL inst_cellmath__63_0_I299 (.Y(N896), .A(N1998), .B(N1834));
NOR2XL inst_cellmath__63_0_I300 (.Y(N898), .A(N1998), .B(N1841));
NOR2XL inst_cellmath__63_0_I301 (.Y(N900), .A(N1998), .B(N1848));
NOR2XL inst_cellmath__63_0_I302 (.Y(N902), .A(N1998), .B(N1855));
NOR2XL inst_cellmath__63_0_I303 (.Y(N904), .A(N1998), .B(N1862));
NOR2XL inst_cellmath__63_0_I304 (.Y(N906), .A(N1998), .B(N1869));
NOR2XL inst_cellmath__63_0_I305 (.Y(N908), .A(N1998), .B(N1876));
NOR2XL inst_cellmath__63_0_I306 (.Y(N910), .A(N1998), .B(N1883));
NOR2XL inst_cellmath__63_0_I307 (.Y(N912), .A(N1998), .B(N1890));
NOR2XL inst_cellmath__63_0_I308 (.Y(N914), .A(N1998), .B(N1897));
NOR2XL inst_cellmath__63_0_I309 (.Y(N916), .A(N1998), .B(N1904));
NOR2XL inst_cellmath__63_0_I310 (.Y(N918), .A(N1998), .B(N1911));
NOR2XL inst_cellmath__63_0_I311 (.Y(N920), .A(N1998), .B(N1918));
NOR2XL inst_cellmath__63_0_I312 (.Y(N922), .A(N1998), .B(N1925));
NOR2XL inst_cellmath__63_0_I313 (.Y(N924), .A(N1998), .B(N1932));
INVXL inst_cellmath__63_0_I1013 (.Y(N2004), .A(inst_cellmath__63_0_in2[11]));
NOR2XL inst_cellmath__63_0_I319 (.Y(N938), .A(N2004), .B(N1813));
NOR2XL inst_cellmath__63_0_I320 (.Y(N940), .A(N2004), .B(N1820));
NOR2XL inst_cellmath__63_0_I321 (.Y(N942), .A(N2004), .B(N1827));
NOR2XL inst_cellmath__63_0_I322 (.Y(N944), .A(N2004), .B(N1834));
NOR2XL inst_cellmath__63_0_I323 (.Y(N946), .A(N2004), .B(N1841));
NOR2XL inst_cellmath__63_0_I324 (.Y(N948), .A(N2004), .B(N1848));
NOR2XL inst_cellmath__63_0_I325 (.Y(N950), .A(N2004), .B(N1855));
NOR2XL inst_cellmath__63_0_I326 (.Y(N952), .A(N2004), .B(N1862));
NOR2XL inst_cellmath__63_0_I327 (.Y(N954), .A(N2004), .B(N1869));
NOR2XL inst_cellmath__63_0_I328 (.Y(N956), .A(N2004), .B(N1876));
NOR2XL inst_cellmath__63_0_I329 (.Y(N958), .A(N2004), .B(N1883));
NOR2XL inst_cellmath__63_0_I330 (.Y(N960), .A(N2004), .B(N1890));
NOR2XL inst_cellmath__63_0_I331 (.Y(N962), .A(N2004), .B(N1897));
NOR2XL inst_cellmath__63_0_I332 (.Y(N964), .A(N2004), .B(N1904));
NOR2XL inst_cellmath__63_0_I333 (.Y(N966), .A(N2004), .B(N1911));
NOR2XL inst_cellmath__63_0_I334 (.Y(N968), .A(N2004), .B(N1918));
NOR2XL inst_cellmath__63_0_I335 (.Y(N970), .A(N2004), .B(N1925));
NOR2XL inst_cellmath__63_0_I336 (.Y(N972), .A(N2004), .B(N1932));
INVXL inst_cellmath__63_0_I1014 (.Y(N2010), .A(inst_cellmath__63_0_in2[12]));
NOR2XL inst_cellmath__63_0_I342 (.Y(N986), .A(N2010), .B(N1813));
NOR2XL inst_cellmath__63_0_I343 (.Y(N988), .A(N2010), .B(N1820));
NOR2XL inst_cellmath__63_0_I344 (.Y(N990), .A(N2010), .B(N1827));
NOR2XL inst_cellmath__63_0_I345 (.Y(N992), .A(N2010), .B(N1834));
NOR2XL inst_cellmath__63_0_I346 (.Y(N994), .A(N2010), .B(N1841));
NOR2XL inst_cellmath__63_0_I347 (.Y(N996), .A(N2010), .B(N1848));
NOR2XL inst_cellmath__63_0_I348 (.Y(N998), .A(N2010), .B(N1855));
NOR2XL inst_cellmath__63_0_I349 (.Y(N1000), .A(N2010), .B(N1862));
NOR2XL inst_cellmath__63_0_I350 (.Y(N1002), .A(N2010), .B(N1869));
NOR2XL inst_cellmath__63_0_I351 (.Y(N1004), .A(N2010), .B(N1876));
NOR2XL inst_cellmath__63_0_I352 (.Y(N1006), .A(N2010), .B(N1883));
NOR2XL inst_cellmath__63_0_I353 (.Y(N1008), .A(N2010), .B(N1890));
NOR2XL inst_cellmath__63_0_I354 (.Y(N1010), .A(N2010), .B(N1897));
NOR2XL inst_cellmath__63_0_I355 (.Y(N1012), .A(N2010), .B(N1904));
NOR2XL inst_cellmath__63_0_I356 (.Y(N1014), .A(N2010), .B(N1911));
NOR2XL inst_cellmath__63_0_I357 (.Y(N1016), .A(N2010), .B(N1918));
NOR2XL inst_cellmath__63_0_I358 (.Y(N1018), .A(N2010), .B(N1925));
NOR2XL inst_cellmath__63_0_I359 (.Y(N1020), .A(N2010), .B(N1932));
INVXL inst_cellmath__63_0_I1015 (.Y(N2016), .A(inst_cellmath__63_0_in2[13]));
NOR2XL inst_cellmath__63_0_I365 (.Y(N1034), .A(N2016), .B(N1813));
NOR2XL inst_cellmath__63_0_I366 (.Y(N1036), .A(N2016), .B(N1820));
NOR2XL inst_cellmath__63_0_I367 (.Y(N1038), .A(N2016), .B(N1827));
NOR2XL inst_cellmath__63_0_I368 (.Y(N1040), .A(N2016), .B(N1834));
NOR2XL inst_cellmath__63_0_I369 (.Y(N1042), .A(N2016), .B(N1841));
NOR2XL inst_cellmath__63_0_I370 (.Y(N1044), .A(N2016), .B(N1848));
NOR2XL inst_cellmath__63_0_I371 (.Y(N1046), .A(N2016), .B(N1855));
NOR2XL inst_cellmath__63_0_I372 (.Y(N1048), .A(N2016), .B(N1862));
NOR2XL inst_cellmath__63_0_I373 (.Y(N1050), .A(N2016), .B(N1869));
NOR2XL inst_cellmath__63_0_I374 (.Y(N1052), .A(N2016), .B(N1876));
NOR2XL inst_cellmath__63_0_I375 (.Y(N1054), .A(N2016), .B(N1883));
NOR2XL inst_cellmath__63_0_I376 (.Y(N1056), .A(N2016), .B(N1890));
NOR2XL inst_cellmath__63_0_I377 (.Y(N1058), .A(N2016), .B(N1897));
NOR2XL inst_cellmath__63_0_I378 (.Y(N1060), .A(N2016), .B(N1904));
NOR2XL inst_cellmath__63_0_I379 (.Y(N1062), .A(N2016), .B(N1911));
NOR2XL inst_cellmath__63_0_I380 (.Y(N1064), .A(N2016), .B(N1918));
NOR2XL inst_cellmath__63_0_I381 (.Y(N1066), .A(N2016), .B(N1925));
NOR2XL inst_cellmath__63_0_I382 (.Y(N1068), .A(N2016), .B(N1932));
INVXL inst_cellmath__63_0_I1016 (.Y(N2022), .A(inst_cellmath__63_0_in2[14]));
NOR2XL inst_cellmath__63_0_I388 (.Y(N1082), .A(N2022), .B(N1813));
NOR2XL inst_cellmath__63_0_I389 (.Y(N1084), .A(N2022), .B(N1820));
NOR2XL inst_cellmath__63_0_I390 (.Y(N1086), .A(N2022), .B(N1827));
NOR2XL inst_cellmath__63_0_I391 (.Y(N1088), .A(N2022), .B(N1834));
NOR2XL inst_cellmath__63_0_I392 (.Y(N1090), .A(N2022), .B(N1841));
NOR2XL inst_cellmath__63_0_I393 (.Y(N1092), .A(N2022), .B(N1848));
NOR2XL inst_cellmath__63_0_I394 (.Y(N1094), .A(N2022), .B(N1855));
NOR2XL inst_cellmath__63_0_I395 (.Y(N1096), .A(N2022), .B(N1862));
NOR2XL inst_cellmath__63_0_I396 (.Y(N1098), .A(N2022), .B(N1869));
NOR2XL inst_cellmath__63_0_I397 (.Y(N1100), .A(N2022), .B(N1876));
NOR2XL inst_cellmath__63_0_I398 (.Y(N1102), .A(N2022), .B(N1883));
NOR2XL inst_cellmath__63_0_I399 (.Y(N1104), .A(N2022), .B(N1890));
NOR2XL inst_cellmath__63_0_I400 (.Y(N1106), .A(N2022), .B(N1897));
NOR2XL inst_cellmath__63_0_I401 (.Y(N1108), .A(N2022), .B(N1904));
NOR2XL inst_cellmath__63_0_I402 (.Y(N1110), .A(N2022), .B(N1911));
NOR2XL inst_cellmath__63_0_I403 (.Y(N1112), .A(N2022), .B(N1918));
NOR2XL inst_cellmath__63_0_I404 (.Y(N1114), .A(N2022), .B(N1925));
NOR2XL inst_cellmath__63_0_I405 (.Y(N1116), .A(N2022), .B(N1932));
NAND2XL inst_cellmath__63_0_I411 (.Y(N1130), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[10]));
NAND2XL inst_cellmath__63_0_I412 (.Y(N1132), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[11]));
NAND2XL inst_cellmath__63_0_I413 (.Y(N1134), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[12]));
NAND2XL inst_cellmath__63_0_I414 (.Y(N1136), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[13]));
NAND2XL inst_cellmath__63_0_I415 (.Y(N1138), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[14]));
NAND2XL inst_cellmath__63_0_I416 (.Y(N1140), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[15]));
NAND2XL inst_cellmath__63_0_I417 (.Y(N1142), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[16]));
NAND2XL inst_cellmath__63_0_I418 (.Y(N1144), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[17]));
NAND2XL inst_cellmath__63_0_I419 (.Y(N1146), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[18]));
NAND2XL inst_cellmath__63_0_I420 (.Y(N1148), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[19]));
NAND2XL inst_cellmath__63_0_I421 (.Y(N1150), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[20]));
NAND2XL inst_cellmath__63_0_I422 (.Y(N1152), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[21]));
NAND2XL inst_cellmath__63_0_I423 (.Y(N1154), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[22]));
NAND2XL inst_cellmath__63_0_I424 (.Y(N1156), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[23]));
NAND2XL inst_cellmath__63_0_I425 (.Y(N1158), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[24]));
NAND2XL inst_cellmath__63_0_I426 (.Y(N1160), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[25]));
NAND2XL inst_cellmath__63_0_I427 (.Y(N1162), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[26]));
NAND2XL inst_cellmath__63_0_I428 (.Y(N1164), .A(inst_cellmath__63_0_in1), .B(inst_cellmath__63_0_in0[27]));
ADDHX1 inst_cellmath__63_0_I446 (.CO(N1185), .S(inst_cellmath__63_0_out0[2]), .A(N414), .B(N506));
ADDHX1 inst_cellmath__63_0_I447 (.CO(N1187), .S(inst_cellmath__63_0_out1[3]), .A(N462), .B(N508));
ADDFX1 inst_cellmath__63_0_I448 (.CO(N1189), .S(inst_cellmath__63_0_out0[3]), .A(N554), .B(N416), .CI(N1185));
ADDHX1 inst_cellmath__63_0_I449 (.CO(N1191), .S(N1190), .A(N510), .B(N556));
ADDFX1 inst_cellmath__63_0_I450 (.CO(N1193), .S(inst_cellmath__63_0_out1[4]), .A(N418), .B(N464), .CI(N602));
ADDFX1 inst_cellmath__63_0_I451 (.CO(inst_cellmath__63_0_out1[5]), .S(inst_cellmath__63_0_out0[4]), .A(N1190), .B(N1187), .CI(N1189));
ADDHX1 inst_cellmath__63_0_I452 (.CO(N1197), .S(N1196), .A(N420), .B(N650));
ADDFX1 inst_cellmath__63_0_I453 (.CO(N1199), .S(N1198), .A(N466), .B(N558), .CI(N512));
ADDFX1 inst_cellmath__63_0_I454 (.CO(N1201), .S(N1200), .A(N1191), .B(N604), .CI(N1196));
ADDFX1 inst_cellmath__63_0_I455 (.CO(inst_cellmath__63_0_out1[6]), .S(inst_cellmath__63_0_out0[5]), .A(N1198), .B(N1193), .CI(N1200));
ADDHX1 inst_cellmath__63_0_I456 (.CO(N1205), .S(N1204), .A(N468), .B(N698));
ADDFX1 inst_cellmath__63_0_I457 (.CO(N1207), .S(N1206), .A(N514), .B(N606), .CI(N560));
ADDFX1 inst_cellmath__63_0_I458 (.CO(N1209), .S(N1208), .A(N652), .B(N422), .CI(N1197));
ADDFX1 inst_cellmath__63_0_I459 (.CO(N1211), .S(N1210), .A(N1204), .B(N1199), .CI(N1206));
ADDFX1 inst_cellmath__63_0_I460 (.CO(inst_cellmath__63_0_out1[7]), .S(inst_cellmath__63_0_out0[6]), .A(N1208), .B(N1201), .CI(N1210));
ADDHX1 inst_cellmath__63_0_I461 (.CO(N1215), .S(N1214), .A(N516), .B(N746));
ADDFX1 inst_cellmath__63_0_I462 (.CO(N1217), .S(N1216), .A(N562), .B(N654), .CI(N424));
ADDFX1 inst_cellmath__63_0_I463 (.CO(N1219), .S(N1218), .A(N470), .B(N608), .CI(N700));
ADDFX1 inst_cellmath__63_0_I464 (.CO(N1221), .S(N1220), .A(N1207), .B(N1205), .CI(N1214));
ADDFX1 inst_cellmath__63_0_I465 (.CO(N1223), .S(N1222), .A(N1209), .B(N1216), .CI(N1218));
ADDFX1 inst_cellmath__63_0_I466 (.CO(inst_cellmath__63_0_out1[8]), .S(inst_cellmath__63_0_out0[7]), .A(N1220), .B(N1211), .CI(N1222));
ADDHX1 inst_cellmath__63_0_I467 (.CO(N1227), .S(N1226), .A(N564), .B(N794));
ADDFX1 inst_cellmath__63_0_I468 (.CO(N1229), .S(N1228), .A(N610), .B(N702), .CI(N426));
ADDFX1 inst_cellmath__63_0_I469 (.CO(N1231), .S(N1230), .A(N472), .B(N656), .CI(N518));
ADDFX1 inst_cellmath__63_0_I470 (.CO(N1233), .S(N1232), .A(N1215), .B(N748), .CI(N1226));
ADDFX1 inst_cellmath__63_0_I471 (.CO(N1235), .S(N1234), .A(N1219), .B(N1217), .CI(N1228));
ADDFX1 inst_cellmath__63_0_I472 (.CO(N1237), .S(N1236), .A(N1221), .B(N1230), .CI(N1232));
ADDFX1 inst_cellmath__63_0_I473 (.CO(inst_cellmath__63_0_out1[9]), .S(inst_cellmath__63_0_out0[8]), .A(N1234), .B(N1223), .CI(N1236));
ADDHX1 inst_cellmath__63_0_I474 (.CO(N1241), .S(N1240), .A(N612), .B(N842));
ADDFX1 inst_cellmath__63_0_I475 (.CO(N1243), .S(N1242), .A(N428), .B(N750), .CI(N474));
ADDFX1 inst_cellmath__63_0_I476 (.CO(N1245), .S(N1244), .A(N658), .B(N704), .CI(N520));
ADDFX1 inst_cellmath__63_0_I477 (.CO(N1247), .S(N1246), .A(N796), .B(N566), .CI(N1227));
ADDFX1 inst_cellmath__63_0_I478 (.CO(N1249), .S(N1248), .A(N1229), .B(N1240), .CI(N1231));
ADDFX1 inst_cellmath__63_0_I479 (.CO(N1251), .S(N1250), .A(N1242), .B(N1244), .CI(N1233));
ADDFX1 inst_cellmath__63_0_I480 (.CO(N1253), .S(N1252), .A(N1235), .B(N1246), .CI(N1248));
ADDFX1 inst_cellmath__63_0_I481 (.CO(inst_cellmath__63_0_out1[10]), .S(inst_cellmath__63_0_out0[9]), .A(N1250), .B(N1237), .CI(N1252));
ADDHX1 inst_cellmath__63_0_I482 (.CO(N1257), .S(N1256), .A(N660), .B(N890));
ADDFX1 inst_cellmath__63_0_I483 (.CO(N1259), .S(N1258), .A(N476), .B(N798), .CI(N522));
ADDFX1 inst_cellmath__63_0_I484 (.CO(N1261), .S(N1260), .A(N706), .B(N430), .CI(N568));
ADDFX1 inst_cellmath__63_0_I485 (.CO(N1263), .S(N1262), .A(N614), .B(N752), .CI(N844));
ADDFX1 inst_cellmath__63_0_I486 (.CO(N1265), .S(N1264), .A(N1256), .B(N1241), .CI(N1243));
ADDFX1 inst_cellmath__63_0_I487 (.CO(N1267), .S(N1266), .A(N1260), .B(N1245), .CI(N1258));
ADDFX1 inst_cellmath__63_0_I488 (.CO(N1269), .S(N1268), .A(N1262), .B(N1247), .CI(N1249));
ADDFX1 inst_cellmath__63_0_I489 (.CO(N1271), .S(N1270), .A(N1251), .B(N1264), .CI(N1266));
ADDFX1 inst_cellmath__63_0_I490 (.CO(inst_cellmath__63_0_out1[11]), .S(inst_cellmath__63_0_out0[10]), .A(N1253), .B(N1268), .CI(N1270));
ADDHX1 inst_cellmath__63_0_I491 (.CO(N1275), .S(N1274), .A(N708), .B(N938));
ADDFX1 inst_cellmath__63_0_I492 (.CO(N1277), .S(N1276), .A(N524), .B(N846), .CI(N570));
ADDFX1 inst_cellmath__63_0_I493 (.CO(N1279), .S(N1278), .A(N754), .B(N478), .CI(N616));
ADDFX1 inst_cellmath__63_0_I494 (.CO(N1281), .S(N1280), .A(N662), .B(N800), .CI(N892));
ADDFX1 inst_cellmath__63_0_I495 (.CO(N1283), .S(N1282), .A(N1257), .B(N432), .CI(N1274));
ADDFX1 inst_cellmath__63_0_I496 (.CO(N1285), .S(N1284), .A(N1259), .B(N1261), .CI(N1263));
ADDFX1 inst_cellmath__63_0_I497 (.CO(N1287), .S(N1286), .A(N1276), .B(N1278), .CI(N1280));
ADDFX1 inst_cellmath__63_0_I498 (.CO(N1289), .S(N1288), .A(N1282), .B(N1265), .CI(N1267));
ADDFX1 inst_cellmath__63_0_I499 (.CO(N1291), .S(N1290), .A(N1269), .B(N1284), .CI(N1286));
ADDFX1 inst_cellmath__63_0_I500 (.CO(inst_cellmath__63_0_out1[12]), .S(inst_cellmath__63_0_out0[11]), .A(N1271), .B(N1288), .CI(N1290));
ADDHX1 inst_cellmath__63_0_I501 (.CO(N1295), .S(N1294), .A(N756), .B(N986));
ADDFX1 inst_cellmath__63_0_I502 (.CO(N1297), .S(N1296), .A(N572), .B(N894), .CI(N618));
ADDFX1 inst_cellmath__63_0_I503 (.CO(N1299), .S(N1298), .A(N802), .B(N526), .CI(N664));
ADDFX1 inst_cellmath__63_0_I504 (.CO(N1301), .S(N1300), .A(N710), .B(N848), .CI(N480));
ADDFX1 inst_cellmath__63_0_I505 (.CO(N1303), .S(N1302), .A(N940), .B(N434), .CI(N1275));
ADDFX1 inst_cellmath__63_0_I506 (.CO(N1305), .S(N1304), .A(N1279), .B(N1294), .CI(N1277));
ADDFX1 inst_cellmath__63_0_I507 (.CO(N1307), .S(N1306), .A(N1298), .B(N1281), .CI(N1296));
ADDFX1 inst_cellmath__63_0_I508 (.CO(N1309), .S(N1308), .A(N1283), .B(N1300), .CI(N1285));
ADDFX1 inst_cellmath__63_0_I509 (.CO(N1311), .S(N1310), .A(N1304), .B(N1302), .CI(N1287));
ADDFX1 inst_cellmath__63_0_I510 (.CO(N1313), .S(N1312), .A(N1289), .B(N1306), .CI(N1308));
ADDFX1 inst_cellmath__63_0_I511 (.CO(inst_cellmath__63_0_out1[13]), .S(inst_cellmath__63_0_out0[12]), .A(N1310), .B(N1291), .CI(N1312));
ADDHX1 inst_cellmath__63_0_I512 (.CO(N1317), .S(N1316), .A(N804), .B(N1034));
ADDFX1 inst_cellmath__63_0_I513 (.CO(N1319), .S(N1318), .A(N436), .B(N942), .CI(N666));
ADDFX1 inst_cellmath__63_0_I514 (.CO(N1321), .S(N1320), .A(N620), .B(N574), .CI(N712));
ADDFX1 inst_cellmath__63_0_I515 (.CO(N1323), .S(N1322), .A(N850), .B(N896), .CI(N758));
ADDFX1 inst_cellmath__63_0_I516 (.CO(N1325), .S(N1324), .A(N988), .B(N482), .CI(N528));
ADDFX1 inst_cellmath__63_0_I517 (.CO(N1327), .S(N1326), .A(N1316), .B(N1295), .CI(N1297));
ADDFX1 inst_cellmath__63_0_I518 (.CO(N1329), .S(N1328), .A(N1301), .B(N1299), .CI(N1320));
ADDFX1 inst_cellmath__63_0_I519 (.CO(N1331), .S(N1330), .A(N1322), .B(N1318), .CI(N1303));
ADDFX1 inst_cellmath__63_0_I520 (.CO(N1333), .S(N1332), .A(N1305), .B(N1324), .CI(N1307));
ADDFX1 inst_cellmath__63_0_I521 (.CO(N1335), .S(N1334), .A(N1328), .B(N1326), .CI(N1309));
ADDFX1 inst_cellmath__63_0_I522 (.CO(N1337), .S(N1336), .A(N1311), .B(N1330), .CI(N1332));
ADDFX1 inst_cellmath__63_0_I523 (.CO(inst_cellmath__63_0_out1[14]), .S(inst_cellmath__63_0_out0[13]), .A(N1313), .B(N1334), .CI(N1336));
ADDHX1 inst_cellmath__63_0_I524 (.CO(N1341), .S(N1340), .A(N438), .B(N484));
ADDFX1 inst_cellmath__63_0_I525 (.CO(N1343), .S(N1342), .A(N990), .B(N852), .CI(N714));
ADDFX1 inst_cellmath__63_0_I526 (.CO(N1345), .S(N1344), .A(N668), .B(N622), .CI(N760));
ADDFX1 inst_cellmath__63_0_I527 (.CO(N1347), .S(N1346), .A(N898), .B(N944), .CI(N806));
ADDFX1 inst_cellmath__63_0_I528 (.CO(N1349), .S(N1348), .A(N1082), .B(N530), .CI(N576));
ADDFX1 inst_cellmath__63_0_I529 (.CO(N1351), .S(N1350), .A(N1317), .B(N1036), .CI(N1340));
ADDFX1 inst_cellmath__63_0_I530 (.CO(N1353), .S(N1352), .A(N1323), .B(N1321), .CI(N1319));
ADDFX1 inst_cellmath__63_0_I531 (.CO(N1355), .S(N1354), .A(N1344), .B(N1325), .CI(N1346));
ADDFX1 inst_cellmath__63_0_I532 (.CO(N1357), .S(N1356), .A(N1348), .B(N1342), .CI(N1327));
ADDFX1 inst_cellmath__63_0_I533 (.CO(N1359), .S(N1358), .A(N1329), .B(N1350), .CI(N1352));
ADDFX1 inst_cellmath__63_0_I534 (.CO(N1361), .S(N1360), .A(N1354), .B(N1331), .CI(N1356));
ADDFX1 inst_cellmath__63_0_I535 (.CO(N1363), .S(N1362), .A(N1358), .B(N1333), .CI(N1335));
ADDFX1 inst_cellmath__63_0_I536 (.CO(inst_cellmath__63_0_out1[15]), .S(inst_cellmath__63_0_out0[14]), .A(N1360), .B(N1337), .CI(N1362));
XNOR2X1 hap1_A_I716 (.Y(N1366), .A(N1130), .B(N440));
OR2XL hap1_A_I717 (.Y(N1367), .A(N1130), .B(N440));
ADDFX1 inst_cellmath__63_0_I538 (.CO(N1371), .S(N1370), .A(N900), .B(N486), .CI(N762));
ADDFX1 inst_cellmath__63_0_I539 (.CO(N1373), .S(N1372), .A(N532), .B(N1038), .CI(N808));
ADDFX1 inst_cellmath__63_0_I540 (.CO(N1375), .S(N1374), .A(N716), .B(N670), .CI(N946));
ADDFX1 inst_cellmath__63_0_I541 (.CO(N1377), .S(N1376), .A(N854), .B(N992), .CI(N624));
ADDFX1 inst_cellmath__63_0_I542 (.CO(N1379), .S(N1378), .A(N1084), .B(N578), .CI(N1341));
ADDFX1 inst_cellmath__63_0_I543 (.CO(N1381), .S(N1380), .A(N1345), .B(N1366), .CI(N1347));
ADDFX1 inst_cellmath__63_0_I544 (.CO(N1383), .S(N1382), .A(N1349), .B(N1343), .CI(N1374));
ADDFX1 inst_cellmath__63_0_I545 (.CO(N1385), .S(N1384), .A(N1370), .B(N1372), .CI(N1376));
ADDFX1 inst_cellmath__63_0_I546 (.CO(N1387), .S(N1386), .A(N1378), .B(N1351), .CI(N1353));
ADDFX1 inst_cellmath__63_0_I547 (.CO(N1389), .S(N1388), .A(N1355), .B(N1380), .CI(N1382));
ADDFX1 inst_cellmath__63_0_I548 (.CO(N1391), .S(N1390), .A(N1384), .B(N1357), .CI(N1359));
ADDFX1 inst_cellmath__63_0_I549 (.CO(N1393), .S(N1392), .A(N1388), .B(N1386), .CI(N1361));
ADDFX1 inst_cellmath__63_0_I550 (.CO(inst_cellmath__63_0_out1[16]), .S(inst_cellmath__63_0_out0[15]), .A(N1363), .B(N1390), .CI(N1392));
ADDFX1 inst_cellmath__63_0_I551 (.CO(N1397), .S(N1396), .A(N1132), .B(N442), .CI(N488));
ADDFX1 inst_cellmath__63_0_I552 (.CO(N1399), .S(N1398), .A(N948), .B(N534), .CI(N810));
ADDFX1 inst_cellmath__63_0_I553 (.CO(N1401), .S(N1400), .A(N580), .B(N1086), .CI(N856));
ADDFX1 inst_cellmath__63_0_I554 (.CO(N1403), .S(N1402), .A(N764), .B(N718), .CI(N994));
ADDFX1 inst_cellmath__63_0_I555 (.CO(N1405), .S(N1404), .A(N902), .B(N1040), .CI(N672));
ADDFX1 inst_cellmath__63_0_I556 (.CO(N1407), .S(N1406), .A(N1367), .B(N626), .CI(N1375));
ADDFX1 inst_cellmath__63_0_I557 (.CO(N1409), .S(N1408), .A(N1371), .B(N1373), .CI(N1396));
ADDFX1 inst_cellmath__63_0_I558 (.CO(N1411), .S(N1410), .A(N1379), .B(N1377), .CI(N1398));
ADDFX1 inst_cellmath__63_0_I559 (.CO(N1413), .S(N1412), .A(N1400), .B(N1402), .CI(N1404));
ADDFX1 inst_cellmath__63_0_I560 (.CO(N1415), .S(N1414), .A(N1383), .B(N1381), .CI(N1406));
ADDFX1 inst_cellmath__63_0_I561 (.CO(N1417), .S(N1416), .A(N1385), .B(N1408), .CI(N1410));
ADDFX1 inst_cellmath__63_0_I562 (.CO(N1419), .S(N1418), .A(N1412), .B(N1387), .CI(N1389));
ADDFX1 inst_cellmath__63_0_I563 (.CO(N1421), .S(N1420), .A(N1391), .B(N1414), .CI(N1416));
ADDFX1 inst_cellmath__63_0_I564 (.CO(inst_cellmath__63_0_out1[17]), .S(inst_cellmath__63_0_out0[16]), .A(N1393), .B(N1418), .CI(N1420));
ADDFX1 inst_cellmath__63_0_I565 (.CO(N1425), .S(N1424), .A(N1134), .B(N444), .CI(N490));
ADDFX1 inst_cellmath__63_0_I566 (.CO(N1427), .S(N1426), .A(N582), .B(N536), .CI(N996));
ADDFX1 inst_cellmath__63_0_I567 (.CO(N1429), .S(N1428), .A(N628), .B(N766), .CI(N858));
ADDFX1 inst_cellmath__63_0_I568 (.CO(N1431), .S(N1430), .A(N812), .B(N1088), .CI(N904));
ADDFX1 inst_cellmath__63_0_I569 (.CO(N1433), .S(N1432), .A(N950), .B(N1042), .CI(N720));
ADDFX1 inst_cellmath__63_0_I570 (.CO(N1435), .S(N1434), .A(N1424), .B(N674), .CI(N1397));
ADDFX1 inst_cellmath__63_0_I571 (.CO(N1437), .S(N1436), .A(N1401), .B(N1403), .CI(N1399));
ADDFX1 inst_cellmath__63_0_I572 (.CO(N1439), .S(N1438), .A(N1426), .B(N1405), .CI(N1430));
ADDFX1 inst_cellmath__63_0_I573 (.CO(N1441), .S(N1440), .A(N1432), .B(N1428), .CI(N1407));
ADDFX1 inst_cellmath__63_0_I574 (.CO(N1443), .S(N1442), .A(N1434), .B(N1409), .CI(N1411));
ADDFX1 inst_cellmath__63_0_I575 (.CO(N1445), .S(N1444), .A(N1413), .B(N1436), .CI(N1438));
ADDFX1 inst_cellmath__63_0_I576 (.CO(N1447), .S(N1446), .A(N1415), .B(N1440), .CI(N1442));
ADDFX1 inst_cellmath__63_0_I577 (.CO(N1449), .S(N1448), .A(N1444), .B(N1417), .CI(N1419));
ADDFX1 inst_cellmath__63_0_I578 (.CO(inst_cellmath__63_0_out1[18]), .S(inst_cellmath__63_0_out0[17]), .A(N1421), .B(N1446), .CI(N1448));
INVXL fap1_A_I718 (.Y(N1803), .A(N1938));
ADDFX1 fap1_A_I719 (.CO(N1453), .S(N1452), .A(N1136), .B(N492), .CI(N1803));
ADDFX1 inst_cellmath__63_0_I580 (.CO(N1457), .S(N1456), .A(N584), .B(N538), .CI(N630));
ADDFX1 inst_cellmath__63_0_I581 (.CO(N1459), .S(N1458), .A(N814), .B(N1044), .CI(N906));
ADDFX1 inst_cellmath__63_0_I582 (.CO(N1461), .S(N1460), .A(N676), .B(N1090), .CI(N722));
ADDFX1 inst_cellmath__63_0_I583 (.CO(N1463), .S(N1462), .A(N952), .B(N860), .CI(N998));
ADDFX1 inst_cellmath__63_0_I584 (.CO(N1465), .S(N1464), .A(N768), .B(N1425), .CI(N1452));
ADDFX1 inst_cellmath__63_0_I585 (.CO(N1467), .S(N1466), .A(N1431), .B(N1427), .CI(N1429));
ADDFX1 inst_cellmath__63_0_I586 (.CO(N1469), .S(N1468), .A(N1433), .B(N1456), .CI(N1458));
ADDFX1 inst_cellmath__63_0_I587 (.CO(N1471), .S(N1470), .A(N1460), .B(N1462), .CI(N1435));
ADDFX1 inst_cellmath__63_0_I588 (.CO(N1473), .S(N1472), .A(N1464), .B(N1437), .CI(N1439));
ADDFX1 inst_cellmath__63_0_I589 (.CO(N1475), .S(N1474), .A(N1441), .B(N1466), .CI(N1468));
ADDFX1 inst_cellmath__63_0_I590 (.CO(N1477), .S(N1476), .A(N1443), .B(N1470), .CI(N1472));
ADDFX1 inst_cellmath__63_0_I591 (.CO(N1479), .S(N1478), .A(N1474), .B(N1445), .CI(N1447));
ADDFX1 inst_cellmath__63_0_I592 (.CO(inst_cellmath__63_0_out1[19]), .S(inst_cellmath__63_0_out0[18]), .A(N1449), .B(N1476), .CI(N1478));
ADDFX1 inst_cellmath__63_0_I593 (.CO(N1483), .S(N1482), .A(N1938), .B(N1944), .CI(N540));
ADDFX1 inst_cellmath__63_0_I594 (.CO(N1485), .S(N1484), .A(N586), .B(N1138), .CI(N1482));
ADDFX1 inst_cellmath__63_0_I595 (.CO(N1487), .S(N1486), .A(N678), .B(N632), .CI(N1092));
ADDFX1 inst_cellmath__63_0_I596 (.CO(N1489), .S(N1488), .A(N1453), .B(N862), .CI(N954));
ADDFX1 inst_cellmath__63_0_I597 (.CO(N1491), .S(N1490), .A(N724), .B(N908), .CI(N770));
ADDFX1 inst_cellmath__63_0_I598 (.CO(N1493), .S(N1492), .A(N1046), .B(N1000), .CI(N816));
ADDFX1 inst_cellmath__63_0_I599 (.CO(N1495), .S(N1494), .A(N1484), .B(N1457), .CI(N1459));
ADDFX1 inst_cellmath__63_0_I600 (.CO(N1497), .S(N1496), .A(N1461), .B(N1463), .CI(N1486));
ADDFX1 inst_cellmath__63_0_I601 (.CO(N1499), .S(N1498), .A(N1465), .B(N1490), .CI(N1492));
ADDFX1 inst_cellmath__63_0_I602 (.CO(N1501), .S(N1500), .A(N1467), .B(N1488), .CI(N1469));
ADDFX1 inst_cellmath__63_0_I603 (.CO(N1503), .S(N1502), .A(N1471), .B(N1494), .CI(N1496));
ADDFX1 inst_cellmath__63_0_I604 (.CO(N1505), .S(N1504), .A(N1473), .B(N1498), .CI(N1500));
ADDFX1 inst_cellmath__63_0_I605 (.CO(N1507), .S(N1506), .A(N1502), .B(N1475), .CI(N1477));
ADDFX1 inst_cellmath__63_0_I606 (.CO(inst_cellmath__63_0_out1[20]), .S(inst_cellmath__63_0_out0[19]), .A(N1479), .B(N1504), .CI(N1506));
ADDFX1 inst_cellmath__63_0_I607 (.CO(N1511), .S(N1510), .A(N588), .B(N1950), .CI(N1483));
ADDFX1 inst_cellmath__63_0_I608 (.CO(N1513), .S(N1512), .A(N634), .B(N1140), .CI(N680));
ADDFX1 inst_cellmath__63_0_I609 (.CO(N1515), .S(N1514), .A(N910), .B(N726), .CI(N1002));
ADDFX1 inst_cellmath__63_0_I610 (.CO(N1517), .S(N1516), .A(N772), .B(N956), .CI(N818));
ADDFX1 inst_cellmath__63_0_I611 (.CO(N1519), .S(N1518), .A(N1094), .B(N1048), .CI(N864));
ADDFX1 inst_cellmath__63_0_I612 (.CO(N1521), .S(N1520), .A(N1510), .B(N1485), .CI(N1487));
ADDFX1 inst_cellmath__63_0_I613 (.CO(N1523), .S(N1522), .A(N1512), .B(N1491), .CI(N1493));
ADDFX1 inst_cellmath__63_0_I614 (.CO(N1525), .S(N1524), .A(N1514), .B(N1489), .CI(N1516));
ADDFX1 inst_cellmath__63_0_I615 (.CO(N1527), .S(N1526), .A(N1495), .B(N1518), .CI(N1497));
ADDFX1 inst_cellmath__63_0_I616 (.CO(N1529), .S(N1528), .A(N1499), .B(N1520), .CI(N1522));
ADDFX1 inst_cellmath__63_0_I617 (.CO(N1531), .S(N1530), .A(N1501), .B(N1524), .CI(N1526));
ADDFX1 inst_cellmath__63_0_I618 (.CO(N1533), .S(N1532), .A(N1528), .B(N1503), .CI(N1505));
ADDFX1 inst_cellmath__63_0_I619 (.CO(inst_cellmath__63_0_out1[21]), .S(inst_cellmath__63_0_out0[20]), .A(N1507), .B(N1530), .CI(N1532));
ADDFX1 inst_cellmath__63_0_I620 (.CO(N1537), .S(N1536), .A(N636), .B(N1956), .CI(N1142));
ADDFX1 inst_cellmath__63_0_I621 (.CO(N1539), .S(N1538), .A(N728), .B(N682), .CI(N774));
ADDFX1 inst_cellmath__63_0_I622 (.CO(N1541), .S(N1540), .A(N958), .B(N1511), .CI(N1050));
ADDFX1 inst_cellmath__63_0_I623 (.CO(N1543), .S(N1542), .A(N820), .B(N1004), .CI(N866));
ADDFX1 inst_cellmath__63_0_I624 (.CO(N1545), .S(N1544), .A(N912), .B(N1096), .CI(N1536));
ADDFX1 inst_cellmath__63_0_I625 (.CO(N1547), .S(N1546), .A(N1515), .B(N1513), .CI(N1517));
ADDFX1 inst_cellmath__63_0_I626 (.CO(N1549), .S(N1548), .A(N1519), .B(N1538), .CI(N1540));
ADDFX1 inst_cellmath__63_0_I627 (.CO(N1551), .S(N1550), .A(N1521), .B(N1542), .CI(N1544));
ADDFX1 inst_cellmath__63_0_I628 (.CO(N1553), .S(N1552), .A(N1546), .B(N1523), .CI(N1525));
ADDFX1 inst_cellmath__63_0_I629 (.CO(N1555), .S(N1554), .A(N1527), .B(N1548), .CI(N1550));
ADDFX1 inst_cellmath__63_0_I630 (.CO(N1557), .S(N1556), .A(N1552), .B(N1529), .CI(N1531));
ADDFX1 inst_cellmath__63_0_I631 (.CO(inst_cellmath__63_0_out1[22]), .S(inst_cellmath__63_0_out0[21]), .A(N1533), .B(N1554), .CI(N1556));
ADDFX1 inst_cellmath__63_0_I632 (.CO(N1561), .S(N1560), .A(N684), .B(N1962), .CI(N1144));
ADDFX1 inst_cellmath__63_0_I633 (.CO(N1563), .S(N1562), .A(N776), .B(N730), .CI(N822));
ADDFX1 inst_cellmath__63_0_I634 (.CO(N1565), .S(N1564), .A(N1537), .B(N1006), .CI(N1098));
ADDFX1 inst_cellmath__63_0_I635 (.CO(N1567), .S(N1566), .A(N868), .B(N1052), .CI(N914));
ADDFX1 inst_cellmath__63_0_I636 (.CO(N1569), .S(N1568), .A(N1560), .B(N960), .CI(N1539));
ADDFX1 inst_cellmath__63_0_I637 (.CO(N1571), .S(N1570), .A(N1543), .B(N1541), .CI(N1562));
ADDFX1 inst_cellmath__63_0_I638 (.CO(N1573), .S(N1572), .A(N1566), .B(N1545), .CI(N1564));
ADDFX1 inst_cellmath__63_0_I639 (.CO(N1575), .S(N1574), .A(N1568), .B(N1547), .CI(N1549));
ADDFX1 inst_cellmath__63_0_I640 (.CO(N1577), .S(N1576), .A(N1551), .B(N1570), .CI(N1572));
ADDFX1 inst_cellmath__63_0_I641 (.CO(N1579), .S(N1578), .A(N1574), .B(N1553), .CI(N1555));
ADDFX1 inst_cellmath__63_0_I642 (.CO(inst_cellmath__63_0_out1[23]), .S(inst_cellmath__63_0_out0[22]), .A(N1557), .B(N1576), .CI(N1578));
ADDFX1 inst_cellmath__63_0_I643 (.CO(N1583), .S(N1582), .A(N732), .B(N1968), .CI(N1146));
ADDFX1 inst_cellmath__63_0_I644 (.CO(N1585), .S(N1584), .A(N824), .B(N778), .CI(N870));
ADDFX1 inst_cellmath__63_0_I645 (.CO(N1587), .S(N1586), .A(N1054), .B(N1561), .CI(N916));
ADDFX1 inst_cellmath__63_0_I646 (.CO(N1589), .S(N1588), .A(N962), .B(N1100), .CI(N1008));
ADDFX1 inst_cellmath__63_0_I647 (.CO(N1591), .S(N1590), .A(N1563), .B(N1582), .CI(N1567));
ADDFX1 inst_cellmath__63_0_I648 (.CO(N1593), .S(N1592), .A(N1584), .B(N1565), .CI(N1586));
ADDFX1 inst_cellmath__63_0_I649 (.CO(N1595), .S(N1594), .A(N1588), .B(N1569), .CI(N1571));
ADDFX1 inst_cellmath__63_0_I650 (.CO(N1597), .S(N1596), .A(N1573), .B(N1590), .CI(N1592));
ADDFX1 inst_cellmath__63_0_I651 (.CO(N1599), .S(N1598), .A(N1594), .B(N1575), .CI(N1577));
ADDFX1 inst_cellmath__63_0_I652 (.CO(inst_cellmath__63_0_out1[24]), .S(inst_cellmath__63_0_out0[23]), .A(N1579), .B(N1596), .CI(N1598));
ADDFX1 inst_cellmath__63_0_I653 (.CO(N1603), .S(N1602), .A(N780), .B(N1974), .CI(N1148));
ADDFX1 inst_cellmath__63_0_I654 (.CO(N1605), .S(N1604), .A(N872), .B(N826), .CI(N918));
ADDFX1 inst_cellmath__63_0_I655 (.CO(N1607), .S(N1606), .A(N1102), .B(N1583), .CI(N964));
ADDFX1 inst_cellmath__63_0_I656 (.CO(N1609), .S(N1608), .A(N1056), .B(N1010), .CI(N1602));
ADDFX1 inst_cellmath__63_0_I657 (.CO(N1611), .S(N1610), .A(N1587), .B(N1585), .CI(N1604));
ADDFX1 inst_cellmath__63_0_I658 (.CO(N1613), .S(N1612), .A(N1606), .B(N1589), .CI(N1608));
ADDFX1 inst_cellmath__63_0_I659 (.CO(N1615), .S(N1614), .A(N1593), .B(N1591), .CI(N1610));
ADDFX1 inst_cellmath__63_0_I660 (.CO(N1617), .S(N1616), .A(N1612), .B(N1595), .CI(N1597));
ADDFX1 inst_cellmath__63_0_I661 (.CO(inst_cellmath__63_0_out1[25]), .S(inst_cellmath__63_0_out0[24]), .A(N1599), .B(N1614), .CI(N1616));
ADDFX1 inst_cellmath__63_0_I662 (.CO(N1621), .S(N1620), .A(N828), .B(N1980), .CI(N1150));
ADDFX1 inst_cellmath__63_0_I663 (.CO(N1623), .S(N1622), .A(N920), .B(N874), .CI(N966));
ADDFX1 inst_cellmath__63_0_I664 (.CO(N1625), .S(N1624), .A(N1012), .B(N1603), .CI(N1058));
ADDFX1 inst_cellmath__63_0_I665 (.CO(N1627), .S(N1626), .A(N1620), .B(N1104), .CI(N1605));
ADDFX1 inst_cellmath__63_0_I666 (.CO(N1629), .S(N1628), .A(N1622), .B(N1607), .CI(N1609));
ADDFX1 inst_cellmath__63_0_I667 (.CO(N1631), .S(N1630), .A(N1626), .B(N1624), .CI(N1611));
ADDFX1 inst_cellmath__63_0_I668 (.CO(N1633), .S(N1632), .A(N1613), .B(N1628), .CI(N1615));
ADDFX1 inst_cellmath__63_0_I669 (.CO(inst_cellmath__63_0_out1[26]), .S(inst_cellmath__63_0_out0[25]), .A(N1617), .B(N1630), .CI(N1632));
ADDFX1 inst_cellmath__63_0_I670 (.CO(N1637), .S(N1636), .A(N876), .B(N1986), .CI(N922));
ADDFX1 inst_cellmath__63_0_I671 (.CO(N1639), .S(N1638), .A(N968), .B(N1152), .CI(N1014));
ADDFX1 inst_cellmath__63_0_I672 (.CO(N1641), .S(N1640), .A(N1060), .B(N1621), .CI(N1106));
ADDFX1 inst_cellmath__63_0_I673 (.CO(N1643), .S(N1642), .A(N1623), .B(N1636), .CI(N1625));
ADDFX1 inst_cellmath__63_0_I674 (.CO(N1645), .S(N1644), .A(N1640), .B(N1638), .CI(N1627));
ADDFX1 inst_cellmath__63_0_I675 (.CO(N1647), .S(N1646), .A(N1642), .B(N1629), .CI(N1644));
ADDFX1 inst_cellmath__63_0_I676 (.CO(inst_cellmath__63_0_out0[27]), .S(inst_cellmath__63_0_out0[26]), .A(N1633), .B(N1631), .CI(N1646));
ADDFX1 inst_cellmath__63_0_I677 (.CO(N1651), .S(N1650), .A(N924), .B(N1992), .CI(N1154));
ADDFX1 inst_cellmath__63_0_I678 (.CO(N1653), .S(N1652), .A(N1016), .B(N970), .CI(N1062));
ADDFX1 inst_cellmath__63_0_I679 (.CO(N1655), .S(N1654), .A(N1637), .B(N1108), .CI(N1650));
ADDFX1 inst_cellmath__63_0_I680 (.CO(N1657), .S(N1656), .A(N1641), .B(N1639), .CI(N1652));
ADDFX1 inst_cellmath__63_0_I681 (.CO(N1659), .S(N1658), .A(N1643), .B(N1654), .CI(N1656));
ADDFX1 inst_cellmath__63_0_I682 (.CO(inst_cellmath__63_0_out0[28]), .S(inst_cellmath__63_0_out1[27]), .A(N1658), .B(N1645), .CI(N1647));
ADDFX1 inst_cellmath__63_0_I683 (.CO(N1663), .S(N1662), .A(N972), .B(N1998), .CI(N1156));
ADDFX1 inst_cellmath__63_0_I684 (.CO(N1665), .S(N1664), .A(N1064), .B(N1018), .CI(N1110));
ADDFX1 inst_cellmath__63_0_I685 (.CO(N1667), .S(N1666), .A(N1662), .B(N1651), .CI(N1653));
ADDFX1 inst_cellmath__63_0_I686 (.CO(N1669), .S(N1668), .A(N1655), .B(N1664), .CI(N1666));
ADDFX1 inst_cellmath__63_0_I687 (.CO(inst_cellmath__63_0_out0[29]), .S(inst_cellmath__63_0_out1[28]), .A(N1668), .B(N1657), .CI(N1659));
ADDFX1 inst_cellmath__63_0_I688 (.CO(N1673), .S(N1672), .A(N1020), .B(N2004), .CI(N1158));
ADDFX1 inst_cellmath__63_0_I689 (.CO(N1675), .S(N1674), .A(N1112), .B(N1066), .CI(N1663));
ADDFX1 inst_cellmath__63_0_I690 (.CO(N1677), .S(N1676), .A(N1665), .B(N1672), .CI(N1674));
ADDFX1 inst_cellmath__63_0_I691 (.CO(inst_cellmath__63_0_out0[30]), .S(inst_cellmath__63_0_out1[29]), .A(N1676), .B(N1667), .CI(N1669));
ADDFX1 inst_cellmath__63_0_I692 (.CO(N1681), .S(N1680), .A(N1068), .B(N2010), .CI(N1160));
ADDFX1 inst_cellmath__63_0_I693 (.CO(N1683), .S(N1682), .A(N1673), .B(N1114), .CI(N1680));
ADDFX1 inst_cellmath__63_0_I694 (.CO(inst_cellmath__63_0_out0[31]), .S(inst_cellmath__63_0_out1[30]), .A(N1682), .B(N1675), .CI(N1677));
ADDFX1 inst_cellmath__63_0_I695 (.CO(N1687), .S(N1686), .A(N1116), .B(N2016), .CI(N1162));
ADDFX1 inst_cellmath__63_0_I696 (.CO(inst_cellmath__63_0_out0[32]), .S(inst_cellmath__63_0_out1[31]), .A(N1686), .B(N1681), .CI(N1683));
ADDFX1 inst_cellmath__63_0_I697 (.CO(inst_cellmath__63_0_out0[33]), .S(inst_cellmath__63_0_out1[32]), .A(N1164), .B(N2022), .CI(N1687));
assign inst_cellmath__63_0_out0[0] = 1'B0;
assign inst_cellmath__63_0_out0[34] = 1'B0;
assign inst_cellmath__63_0_out0[35] = 1'B0;
assign inst_cellmath__63_0_out0[36] = 1'B0;
assign inst_cellmath__63_0_out0[37] = 1'B0;
assign inst_cellmath__63_0_out0[38] = 1'B0;
assign inst_cellmath__63_0_out0[39] = 1'B0;
assign inst_cellmath__63_0_out1[33] = inst_cellmath__63_0_in1;
assign inst_cellmath__63_0_out1[34] = 1'B1;
assign inst_cellmath__63_0_out1[35] = 1'B1;
assign inst_cellmath__63_0_out1[36] = 1'B1;
assign inst_cellmath__63_0_out1[37] = 1'B1;
assign inst_cellmath__63_0_out1[38] = 1'B1;
assign inst_cellmath__63_0_out1[39] = 1'B1;
endmodule

module cynw_cm_float_rcp_inst_cellmath__64_0_bdw1412651405_bdw (
	inst_cellmath__64_0_out0,
	inst_cellmath__64_0_in0,
	inst_cellmath__64_0_in1,
	inst_cellmath__64_0_in2,
	inst_cellmath__64_0_in3,
	inst_cellmath__64_0_in4
	); /* architecture "gate_level" */ 
output [39:0] inst_cellmath__64_0_out0;
input [52:28] inst_cellmath__64_0_in0;
input [39:0] inst_cellmath__64_0_in1,
	inst_cellmath__64_0_in2,
	inst_cellmath__64_0_in3,
	inst_cellmath__64_0_in4;
wire N1509,N1510,N1511,N1512,N1515,N1516,N1517 
	,N1518,N1519,N1520,N1521,N1522,N1523,N1524,N1525 
	,N1526,N1527,N1528,N1529,N1530,N1531,N1532,N1533 
	,N1534,N1535,N1536,N1537,N1538,N1539,N1540,N1541 
	,N1542,N1543,N1544,N1545,N1546,N1547,N1548,N1549 
	,N1550,N1551,N1552,N1553,N1554,N1555,N1556,N1557 
	,N1558,N1559,N1560,N1561,N1562,N1563,N1564,N1565 
	,N1566,N1567,N1568,N1569,N1570,N1571,N1572,N1573 
	,N1574,N1575,N1576,N1577,N1578,N1579,N1580,N1581 
	,N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589 
	,N1590,N1591,N1592,N1593,N1594,N1595,N1596,N1597 
	,N1598,N1599,N1600,N1601,N1602,N1603,N1604,N1605 
	,N1606,N1607,N1609,N1610,N1611,N1612,N1613,N1614 
	,N1615,N1616,N1617,N1618,N1619,N1620,N1621,N1622 
	,N1623,N1624,N1625,N1626,N1627,N1628,N1629,N1630 
	,N1631,N1632,N1633,N1634,N1635,N1636,N1637,N1638 
	,N1639,N1640,N1641,N1642,N1643,N1644,N1645,N1646 
	,N1647,N1648,N1649,N1650,N1651,N1652,N1653,N1654 
	,N1655,N1656,N1657,N1658,N1659,N1660,N1661,N1662 
	,N1663,N1664,N1665,N1666,N1667,N1668,N1669,N1670 
	,N1671,N1672,N1673,N1674,N1675,N1676,N1677,N1678 
	,N1679,N1680,N1681,N1682,N1683,N1684,N1685,N1686 
	,N1687,N1688,N1689,N1690,N1691,N1692,N1693,N1694 
	,N1695,N1696,N1697,N1698,N1699,N1700,N1701,N1702 
	,N1703,N1704,N1705,N1706,N1707,N1708,N1709,N1710 
	,N1711,N1712,N1713,N1714,N1715,N1716,N1717,N1718 
	,N1719,N1720,N1721,N1722,N1723,N1724,N1725,N1726 
	,N1727,N1728,N1729,N1730,N1731,N1732,N1733,N1734 
	,N1735,N1736,N1737,N1738,N1739,N1740,N1741,N1742 
	,N1743,N1744,N1745,N1746,N1747,N1748,N1749,N1750 
	,N1751,N1752,N1753,N1754,N1755,N1756,N1759,N1767 
	,N1775,N1787,N1799,N1815,N1831,N1851,N1871,N1895 
	,N1919,N1947,N1975,N2014,N2017,N2020,N2023,N2026 
	,N2029,N2032,N2035,N2038,N2041,N2044,N2047,N2050 
	,N2053,N2070,N2072,N2073,N2075,N2077,N2079,N2081 
	,N2083,N2085,N2087,N2089,N2091,N2093,N2095,N2097 
	,N2099,N2101,N2103,N2105,N2107,N2109,N2111,N2113 
	,N2115,N2117,N2119,N2121,N2124,N2132,N2140,N2152 
	,N2164,N2180,N2196,N2216,N2236,N2260,N2284,N2312 
	,N2340,N2372,N2404,N2440,N2476,N2516,N2556,N2600 
	,N2644,N2692,N2740,N3161,N3167,N3180,N3193,N3206 
	,N3219,N3232,N3245,N3258,N3271,N3284,N3297,N3310 
	,N3323,N3336,N3349,N3362,N3375,N3388,N3401,N3414 
	,N3427,N3440,N3453,N3466,N3479,N3492,N3505,N3518 
	,N3531,N3544,N3557,N3570,N3583,N3596,N3609,N3622 
	,N3635,N3648,N3721,N3722,N3728,N3729,N3743,N3744 
	,N3762,N3763,N3785,N3786,N3812,N3813,N3843,N3844 
	,N4195;
ADDHX1 inst_cellmath__64_0_I412 (.CO(N1510), .S(N1509), .A(inst_cellmath__64_0_in0[28]), .B(inst_cellmath__64_0_in2[15]));
XNOR2X1 hap1_A_I1749 (.Y(N1511), .A(inst_cellmath__64_0_in0[29]), .B(inst_cellmath__64_0_in2[16]));
OR2XL hap1_A_I1750 (.Y(N1512), .A(inst_cellmath__64_0_in0[29]), .B(inst_cellmath__64_0_in2[16]));
ADDHX1 inst_cellmath__64_0_I414 (.CO(N1516), .S(N1515), .A(inst_cellmath__64_0_in1[16]), .B(inst_cellmath__64_0_in4[16]));
ADDFX1 inst_cellmath__64_0_I415 (.CO(N1518), .S(N1517), .A(inst_cellmath__64_0_in2[17]), .B(inst_cellmath__64_0_in0[30]), .CI(inst_cellmath__64_0_in1[17]));
ADDHX1 inst_cellmath__64_0_I416 (.CO(N1520), .S(N1519), .A(inst_cellmath__64_0_in4[17]), .B(inst_cellmath__64_0_in3[17]));
ADDFX1 inst_cellmath__64_0_I417 (.CO(N1522), .S(N1521), .A(inst_cellmath__64_0_in2[18]), .B(inst_cellmath__64_0_in0[31]), .CI(inst_cellmath__64_0_in1[18]));
ADDHX1 inst_cellmath__64_0_I418 (.CO(N1524), .S(N1523), .A(inst_cellmath__64_0_in4[18]), .B(inst_cellmath__64_0_in3[18]));
ADDFX1 inst_cellmath__64_0_I419 (.CO(N1526), .S(N1525), .A(inst_cellmath__64_0_in2[19]), .B(inst_cellmath__64_0_in0[32]), .CI(inst_cellmath__64_0_in1[19]));
ADDHX1 inst_cellmath__64_0_I420 (.CO(N1528), .S(N1527), .A(inst_cellmath__64_0_in4[19]), .B(inst_cellmath__64_0_in3[19]));
ADDFX1 inst_cellmath__64_0_I421 (.CO(N1530), .S(N1529), .A(inst_cellmath__64_0_in2[20]), .B(inst_cellmath__64_0_in0[33]), .CI(inst_cellmath__64_0_in1[20]));
ADDHX1 inst_cellmath__64_0_I422 (.CO(N1532), .S(N1531), .A(inst_cellmath__64_0_in4[20]), .B(inst_cellmath__64_0_in3[20]));
ADDFX1 inst_cellmath__64_0_I423 (.CO(N1534), .S(N1533), .A(inst_cellmath__64_0_in2[21]), .B(inst_cellmath__64_0_in0[34]), .CI(inst_cellmath__64_0_in1[21]));
ADDHX1 inst_cellmath__64_0_I424 (.CO(N1536), .S(N1535), .A(inst_cellmath__64_0_in4[21]), .B(inst_cellmath__64_0_in3[21]));
ADDFX1 inst_cellmath__64_0_I425 (.CO(N1538), .S(N1537), .A(inst_cellmath__64_0_in2[22]), .B(inst_cellmath__64_0_in0[35]), .CI(inst_cellmath__64_0_in4[22]));
ADDHX1 inst_cellmath__64_0_I426 (.CO(N1540), .S(N1539), .A(inst_cellmath__64_0_in1[22]), .B(inst_cellmath__64_0_in3[22]));
ADDFX1 inst_cellmath__64_0_I427 (.CO(N1542), .S(N1541), .A(inst_cellmath__64_0_in4[23]), .B(inst_cellmath__64_0_in0[36]), .CI(inst_cellmath__64_0_in3[23]));
ADDHX1 inst_cellmath__64_0_I428 (.CO(N1544), .S(N1543), .A(inst_cellmath__64_0_in2[23]), .B(inst_cellmath__64_0_in1[23]));
ADDFX1 inst_cellmath__64_0_I429 (.CO(N1546), .S(N1545), .A(inst_cellmath__64_0_in4[24]), .B(inst_cellmath__64_0_in0[37]), .CI(inst_cellmath__64_0_in3[24]));
ADDHX1 inst_cellmath__64_0_I430 (.CO(N1548), .S(N1547), .A(inst_cellmath__64_0_in2[24]), .B(inst_cellmath__64_0_in1[24]));
ADDFX1 inst_cellmath__64_0_I431 (.CO(N1550), .S(N1549), .A(inst_cellmath__64_0_in3[25]), .B(inst_cellmath__64_0_in4[25]), .CI(inst_cellmath__64_0_in0[38]));
ADDHX1 inst_cellmath__64_0_I432 (.CO(N1552), .S(N1551), .A(inst_cellmath__64_0_in2[25]), .B(inst_cellmath__64_0_in1[25]));
ADDFX1 inst_cellmath__64_0_I433 (.CO(N1554), .S(N1553), .A(inst_cellmath__64_0_in3[26]), .B(inst_cellmath__64_0_in4[26]), .CI(inst_cellmath__64_0_in0[39]));
ADDHX1 inst_cellmath__64_0_I434 (.CO(N1556), .S(N1555), .A(inst_cellmath__64_0_in2[26]), .B(inst_cellmath__64_0_in1[26]));
ADDFX1 inst_cellmath__64_0_I435 (.CO(N1558), .S(N1557), .A(inst_cellmath__64_0_in3[27]), .B(inst_cellmath__64_0_in4[27]), .CI(inst_cellmath__64_0_in0[40]));
ADDHX1 inst_cellmath__64_0_I436 (.CO(N1560), .S(N1559), .A(inst_cellmath__64_0_in2[27]), .B(inst_cellmath__64_0_in1[27]));
ADDFX1 inst_cellmath__64_0_I437 (.CO(N1562), .S(N1561), .A(inst_cellmath__64_0_in3[28]), .B(inst_cellmath__64_0_in4[28]), .CI(inst_cellmath__64_0_in0[41]));
ADDHX1 inst_cellmath__64_0_I438 (.CO(N1564), .S(N1563), .A(inst_cellmath__64_0_in2[28]), .B(inst_cellmath__64_0_in1[28]));
ADDFX1 inst_cellmath__64_0_I439 (.CO(N1566), .S(N1565), .A(inst_cellmath__64_0_in3[29]), .B(inst_cellmath__64_0_in4[29]), .CI(inst_cellmath__64_0_in0[42]));
ADDHX1 inst_cellmath__64_0_I440 (.CO(N1568), .S(N1567), .A(inst_cellmath__64_0_in2[29]), .B(inst_cellmath__64_0_in1[29]));
ADDFX1 inst_cellmath__64_0_I441 (.CO(N1570), .S(N1569), .A(inst_cellmath__64_0_in3[30]), .B(inst_cellmath__64_0_in4[30]), .CI(inst_cellmath__64_0_in0[43]));
ADDHX1 inst_cellmath__64_0_I442 (.CO(N1572), .S(N1571), .A(inst_cellmath__64_0_in2[30]), .B(inst_cellmath__64_0_in1[30]));
ADDFX1 inst_cellmath__64_0_I443 (.CO(N1574), .S(N1573), .A(inst_cellmath__64_0_in3[31]), .B(inst_cellmath__64_0_in4[31]), .CI(inst_cellmath__64_0_in0[44]));
ADDHX1 inst_cellmath__64_0_I444 (.CO(N1576), .S(N1575), .A(inst_cellmath__64_0_in2[31]), .B(inst_cellmath__64_0_in1[31]));
ADDFX1 inst_cellmath__64_0_I445 (.CO(N1578), .S(N1577), .A(inst_cellmath__64_0_in3[32]), .B(inst_cellmath__64_0_in4[32]), .CI(inst_cellmath__64_0_in0[45]));
ADDHX1 inst_cellmath__64_0_I446 (.CO(N1580), .S(N1579), .A(inst_cellmath__64_0_in2[32]), .B(inst_cellmath__64_0_in1[32]));
ADDFX1 inst_cellmath__64_0_I447 (.CO(N1582), .S(N1581), .A(inst_cellmath__64_0_in3[33]), .B(inst_cellmath__64_0_in4[33]), .CI(inst_cellmath__64_0_in2[33]));
ADDHX1 inst_cellmath__64_0_I448 (.CO(N1584), .S(N1583), .A(inst_cellmath__64_0_in0[46]), .B(inst_cellmath__64_0_in1[33]));
ADDFX1 inst_cellmath__64_0_I449 (.CO(N1586), .S(N1585), .A(inst_cellmath__64_0_in1[34]), .B(inst_cellmath__64_0_in2[34]), .CI(inst_cellmath__64_0_in4[34]));
ADDHX1 inst_cellmath__64_0_I450 (.CO(N1588), .S(N1587), .A(inst_cellmath__64_0_in3[34]), .B(inst_cellmath__64_0_in0[47]));
ADDFX1 inst_cellmath__64_0_I451 (.CO(N1590), .S(N1589), .A(inst_cellmath__64_0_in1[35]), .B(inst_cellmath__64_0_in2[35]), .CI(inst_cellmath__64_0_in4[35]));
ADDHX1 inst_cellmath__64_0_I452 (.CO(N1592), .S(N1591), .A(inst_cellmath__64_0_in3[35]), .B(inst_cellmath__64_0_in0[48]));
ADDFX1 inst_cellmath__64_0_I453 (.CO(N1594), .S(N1593), .A(inst_cellmath__64_0_in1[36]), .B(inst_cellmath__64_0_in2[36]), .CI(inst_cellmath__64_0_in4[36]));
ADDHX1 inst_cellmath__64_0_I454 (.CO(N1596), .S(N1595), .A(inst_cellmath__64_0_in3[36]), .B(inst_cellmath__64_0_in0[49]));
ADDFX1 inst_cellmath__64_0_I455 (.CO(N1598), .S(N1597), .A(inst_cellmath__64_0_in1[37]), .B(inst_cellmath__64_0_in2[37]), .CI(inst_cellmath__64_0_in4[37]));
ADDHX1 inst_cellmath__64_0_I456 (.CO(N1600), .S(N1599), .A(inst_cellmath__64_0_in3[37]), .B(inst_cellmath__64_0_in0[50]));
ADDFX1 inst_cellmath__64_0_I457 (.CO(N1602), .S(N1601), .A(inst_cellmath__64_0_in1[38]), .B(inst_cellmath__64_0_in2[38]), .CI(inst_cellmath__64_0_in4[38]));
ADDHX1 inst_cellmath__64_0_I458 (.CO(N1604), .S(N1603), .A(inst_cellmath__64_0_in3[38]), .B(inst_cellmath__64_0_in0[51]));
ADDFX1 inst_cellmath__64_0_I459 (.CO(N1606), .S(N1605), .A(inst_cellmath__64_0_in1[39]), .B(inst_cellmath__64_0_in2[39]), .CI(inst_cellmath__64_0_in4[39]));
XOR2XL inst_cellmath__64_0_I460 (.Y(N1607), .A(inst_cellmath__64_0_in3[39]), .B(inst_cellmath__64_0_in0[52]));
ADDFX1 inst_cellmath__64_0_I461 (.CO(N1610), .S(N1609), .A(inst_cellmath__64_0_in4[0]), .B(inst_cellmath__64_0_in1[0]), .CI(inst_cellmath__64_0_in3[0]));
ADDHX1 arith_dha_A_I1751 (.CO(N1612), .S(N3161), .A(inst_cellmath__64_0_in4[1]), .B(inst_cellmath__64_0_in3[1]));
ADDFX1 arith_dha_A_I1752 (.CO(N1613), .S(N1611), .A(N3161), .B(inst_cellmath__64_0_in2[1]), .CI(inst_cellmath__64_0_in1[1]));
ADDFX1 arith_dfa_A_I1753 (.CO(N1616), .S(N3167), .A(inst_cellmath__64_0_in3[2]), .B(inst_cellmath__64_0_in4[2]), .CI(inst_cellmath__64_0_in2[2]));
ADDFX1 arith_dfa_A_I1754 (.CO(N1615), .S(N1614), .A(N1612), .B(inst_cellmath__64_0_in1[2]), .CI(N3167));
ADDFX1 arith_dfa_A_I1755 (.CO(N1619), .S(N3180), .A(inst_cellmath__64_0_in3[3]), .B(inst_cellmath__64_0_in4[3]), .CI(inst_cellmath__64_0_in2[3]));
ADDFX1 arith_dfa_A_I1756 (.CO(N1618), .S(N1617), .A(N1616), .B(inst_cellmath__64_0_in1[3]), .CI(N3180));
ADDFX1 arith_dfa_A_I1757 (.CO(N1622), .S(N3193), .A(inst_cellmath__64_0_in2[4]), .B(inst_cellmath__64_0_in3[4]), .CI(inst_cellmath__64_0_in4[4]));
ADDFX1 arith_dfa_A_I1758 (.CO(N1621), .S(N1620), .A(inst_cellmath__64_0_in1[4]), .B(N1619), .CI(N3193));
ADDFX1 arith_dfa_A_I1759 (.CO(N1625), .S(N3206), .A(inst_cellmath__64_0_in3[5]), .B(inst_cellmath__64_0_in2[5]), .CI(inst_cellmath__64_0_in4[5]));
ADDFX1 arith_dfa_A_I1760 (.CO(N1624), .S(N1623), .A(N1622), .B(inst_cellmath__64_0_in1[5]), .CI(N3206));
ADDFX1 arith_dfa_A_I1761 (.CO(N1628), .S(N3219), .A(inst_cellmath__64_0_in2[6]), .B(inst_cellmath__64_0_in4[6]), .CI(inst_cellmath__64_0_in3[6]));
ADDFX1 arith_dfa_A_I1762 (.CO(N1627), .S(N1626), .A(N1625), .B(inst_cellmath__64_0_in1[6]), .CI(N3219));
ADDFX1 arith_dfa_A_I1763 (.CO(N1631), .S(N3232), .A(inst_cellmath__64_0_in2[7]), .B(inst_cellmath__64_0_in4[7]), .CI(inst_cellmath__64_0_in1[7]));
ADDFX1 arith_dfa_A_I1764 (.CO(N1630), .S(N1629), .A(inst_cellmath__64_0_in3[7]), .B(N1628), .CI(N3232));
ADDFX1 arith_dfa_A_I1765 (.CO(N1634), .S(N3245), .A(inst_cellmath__64_0_in4[8]), .B(inst_cellmath__64_0_in2[8]), .CI(inst_cellmath__64_0_in1[8]));
ADDFX1 arith_dfa_A_I1766 (.CO(N1633), .S(N1632), .A(N1631), .B(inst_cellmath__64_0_in3[8]), .CI(N3245));
ADDFX1 arith_dfa_A_I1767 (.CO(N1637), .S(N3258), .A(inst_cellmath__64_0_in1[9]), .B(inst_cellmath__64_0_in2[9]), .CI(inst_cellmath__64_0_in4[9]));
ADDFX1 arith_dfa_A_I1768 (.CO(N1636), .S(N1635), .A(N1634), .B(inst_cellmath__64_0_in3[9]), .CI(N3258));
ADDFX1 arith_dfa_A_I1769 (.CO(N1640), .S(N3271), .A(inst_cellmath__64_0_in1[10]), .B(inst_cellmath__64_0_in2[10]), .CI(inst_cellmath__64_0_in4[10]));
ADDFX1 arith_dfa_A_I1770 (.CO(N1639), .S(N1638), .A(N1637), .B(inst_cellmath__64_0_in3[10]), .CI(N3271));
ADDFX1 arith_dfa_A_I1771 (.CO(N1643), .S(N3284), .A(inst_cellmath__64_0_in1[11]), .B(inst_cellmath__64_0_in2[11]), .CI(inst_cellmath__64_0_in4[11]));
ADDFX1 arith_dfa_A_I1772 (.CO(N1642), .S(N1641), .A(N1640), .B(inst_cellmath__64_0_in3[11]), .CI(N3284));
ADDFX1 arith_dfa_A_I1773 (.CO(N1646), .S(N3297), .A(inst_cellmath__64_0_in1[12]), .B(inst_cellmath__64_0_in2[12]), .CI(inst_cellmath__64_0_in4[12]));
ADDFX1 arith_dfa_A_I1774 (.CO(N1645), .S(N1644), .A(N3297), .B(N1643), .CI(inst_cellmath__64_0_in3[12]));
ADDFX1 arith_dfa_A_I1775 (.CO(N1649), .S(N3310), .A(inst_cellmath__64_0_in1[13]), .B(inst_cellmath__64_0_in2[13]), .CI(inst_cellmath__64_0_in4[13]));
ADDFX1 arith_dfa_A_I1776 (.CO(N1648), .S(N1647), .A(N1646), .B(inst_cellmath__64_0_in3[13]), .CI(N3310));
ADDFX1 arith_dfa_A_I1777 (.CO(N1652), .S(N3323), .A(inst_cellmath__64_0_in1[14]), .B(inst_cellmath__64_0_in2[14]), .CI(inst_cellmath__64_0_in4[14]));
ADDFX1 arith_dfa_A_I1778 (.CO(N1651), .S(N1650), .A(N1649), .B(inst_cellmath__64_0_in3[14]), .CI(N3323));
ADDFX1 arith_dfa_A_I1779 (.CO(N1655), .S(N3336), .A(inst_cellmath__64_0_in1[15]), .B(N1509), .CI(inst_cellmath__64_0_in4[15]));
ADDFX1 arith_dfa_A_I1780 (.CO(N1654), .S(N1653), .A(N1652), .B(inst_cellmath__64_0_in3[15]), .CI(N3336));
ADDFX1 arith_dfa_A_I1781 (.CO(N1658), .S(N3349), .A(N1511), .B(N1510), .CI(inst_cellmath__64_0_in3[16]));
ADDFX1 arith_dfa_A_I1782 (.CO(N1657), .S(N1656), .A(N1655), .B(N1515), .CI(N3349));
ADDFX1 arith_dfa_A_I1783 (.CO(N1661), .S(N3362), .A(N1517), .B(N1512), .CI(N1516));
ADDFX1 arith_dfa_A_I1784 (.CO(N1660), .S(N1659), .A(N1658), .B(N1519), .CI(N3362));
ADDFX1 arith_dfa_A_I1785 (.CO(N1664), .S(N3375), .A(N1521), .B(N1518), .CI(N1523));
ADDFX1 arith_dfa_A_I1786 (.CO(N1663), .S(N1662), .A(N1661), .B(N1520), .CI(N3375));
ADDFX1 arith_dfa_A_I1787 (.CO(N1667), .S(N3388), .A(N1525), .B(N1522), .CI(N1527));
ADDFX1 arith_dfa_A_I1788 (.CO(N1666), .S(N1665), .A(N1664), .B(N1524), .CI(N3388));
ADDFX1 arith_dfa_A_I1789 (.CO(N1670), .S(N3401), .A(N1529), .B(N1526), .CI(N1528));
ADDFX1 arith_dfa_A_I1790 (.CO(N1669), .S(N1668), .A(N1667), .B(N1531), .CI(N3401));
ADDFX1 arith_dfa_A_I1791 (.CO(N1673), .S(N3414), .A(N1533), .B(N1530), .CI(N1535));
ADDFX1 arith_dfa_A_I1792 (.CO(N1672), .S(N1671), .A(N1670), .B(N1532), .CI(N3414));
ADDFX1 arith_dfa_A_I1793 (.CO(N1676), .S(N3427), .A(N1539), .B(N1534), .CI(N1537));
ADDFX1 arith_dfa_A_I1794 (.CO(N1675), .S(N1674), .A(N1673), .B(N1536), .CI(N3427));
ADDFX1 arith_dfa_A_I1795 (.CO(N1679), .S(N3440), .A(N1541), .B(N1543), .CI(N1540));
ADDFX1 arith_dfa_A_I1796 (.CO(N1678), .S(N1677), .A(N1676), .B(N1538), .CI(N3440));
ADDFX1 arith_dfa_A_I1797 (.CO(N1682), .S(N3453), .A(N1547), .B(N1545), .CI(N1544));
ADDFX1 arith_dfa_A_I1798 (.CO(N1681), .S(N1680), .A(N1679), .B(N1542), .CI(N3453));
ADDFX1 arith_dfa_A_I1799 (.CO(N1685), .S(N3466), .A(N1546), .B(N1549), .CI(N1548));
ADDFX1 arith_dfa_A_I1800 (.CO(N1684), .S(N1683), .A(N1682), .B(N1551), .CI(N3466));
ADDFX1 arith_dfa_A_I1801 (.CO(N1688), .S(N3479), .A(N1553), .B(N1550), .CI(N1555));
ADDFX1 arith_dfa_A_I1802 (.CO(N1687), .S(N1686), .A(N1685), .B(N1552), .CI(N3479));
ADDFX1 arith_dfa_A_I1803 (.CO(N1691), .S(N3492), .A(N1557), .B(N1554), .CI(N1559));
ADDFX1 arith_dfa_A_I1804 (.CO(N1690), .S(N1689), .A(N1688), .B(N1556), .CI(N3492));
ADDFX1 arith_dfa_A_I1805 (.CO(N1694), .S(N3505), .A(N1561), .B(N1558), .CI(N1563));
ADDFX1 arith_dfa_A_I1806 (.CO(N1693), .S(N1692), .A(N1691), .B(N1560), .CI(N3505));
ADDFX1 arith_dfa_A_I1807 (.CO(N1697), .S(N3518), .A(N1565), .B(N1562), .CI(N1567));
ADDFX1 arith_dfa_A_I1808 (.CO(N1696), .S(N1695), .A(N1694), .B(N1564), .CI(N3518));
ADDFX1 arith_dfa_A_I1809 (.CO(N1700), .S(N3531), .A(N1569), .B(N1566), .CI(N1571));
ADDFX1 arith_dfa_A_I1810 (.CO(N1699), .S(N1698), .A(N1697), .B(N1568), .CI(N3531));
ADDFX1 arith_dfa_A_I1811 (.CO(N1703), .S(N3544), .A(N1573), .B(N1570), .CI(N1575));
ADDFX1 arith_dfa_A_I1812 (.CO(N1702), .S(N1701), .A(N1700), .B(N1572), .CI(N3544));
ADDFX1 arith_dfa_A_I1813 (.CO(N1706), .S(N3557), .A(N1577), .B(N1574), .CI(N1579));
ADDFX1 arith_dfa_A_I1814 (.CO(N1705), .S(N1704), .A(N1703), .B(N1576), .CI(N3557));
ADDFX1 arith_dfa_A_I1815 (.CO(N1709), .S(N3570), .A(N1578), .B(N1581), .CI(N1583));
ADDFX1 arith_dfa_A_I1816 (.CO(N1708), .S(N1707), .A(N1706), .B(N1580), .CI(N3570));
ADDFX1 arith_dfa_A_I1817 (.CO(N1712), .S(N3583), .A(N1582), .B(N1585), .CI(N1587));
ADDFX1 arith_dfa_A_I1818 (.CO(N1711), .S(N1710), .A(N1709), .B(N1584), .CI(N3583));
ADDFX1 arith_dfa_A_I1819 (.CO(N1715), .S(N3596), .A(N1589), .B(N1586), .CI(N1588));
ADDFX1 arith_dfa_A_I1820 (.CO(N1714), .S(N1713), .A(N1712), .B(N1591), .CI(N3596));
ADDFX1 arith_dfa_A_I1821 (.CO(N1718), .S(N3609), .A(N1593), .B(N1590), .CI(N1595));
ADDFX1 arith_dfa_A_I1822 (.CO(N1717), .S(N1716), .A(N1715), .B(N1592), .CI(N3609));
ADDFX1 arith_dfa_A_I1823 (.CO(N1721), .S(N3622), .A(N1597), .B(N1594), .CI(N1599));
ADDFX1 arith_dfa_A_I1824 (.CO(N1720), .S(N1719), .A(N1718), .B(N1596), .CI(N3622));
ADDFX1 arith_dfa_A_I1825 (.CO(N1724), .S(N3635), .A(N1601), .B(N1598), .CI(N1600));
ADDFX1 arith_dfa_A_I1826 (.CO(N1723), .S(N1722), .A(N1721), .B(N1603), .CI(N3635));
ADDFX1 arith_dfa_A_I1827 (.CO(N1727), .S(N3648), .A(N1605), .B(N1602), .CI(N1607));
ADDFX1 arith_dfa_A_I1828 (.CO(N1726), .S(N1725), .A(N1724), .B(N1604), .CI(N3648));
NAND2XL inst_cellmath__64_0_I501 (.Y(N1728), .A(N1609), .B(inst_cellmath__64_0_in2[0]));
NOR2XL inst_cellmath__64_0_I502 (.Y(N1729), .A(N1610), .B(N1611));
NAND2XL inst_cellmath__64_0_I503 (.Y(N1730), .A(N1610), .B(N1611));
NOR2XL inst_cellmath__64_0_I504 (.Y(N1731), .A(N1613), .B(N1614));
NAND2XL inst_cellmath__64_0_I505 (.Y(N1732), .A(N1613), .B(N1614));
NOR2XL inst_cellmath__64_0_I506 (.Y(N1733), .A(N1615), .B(N1617));
NAND2XL inst_cellmath__64_0_I507 (.Y(N1734), .A(N1615), .B(N1617));
NOR2XL inst_cellmath__64_0_I508 (.Y(N1735), .A(N1618), .B(N1620));
NAND2XL inst_cellmath__64_0_I509 (.Y(N1736), .A(N1618), .B(N1620));
NOR2XL inst_cellmath__64_0_I510 (.Y(N1737), .A(N1621), .B(N1623));
NAND2XL inst_cellmath__64_0_I511 (.Y(N1738), .A(N1621), .B(N1623));
NOR2XL inst_cellmath__64_0_I512 (.Y(N1739), .A(N1624), .B(N1626));
NAND2XL inst_cellmath__64_0_I513 (.Y(N1740), .A(N1624), .B(N1626));
NOR2XL inst_cellmath__64_0_I514 (.Y(N1741), .A(N1627), .B(N1629));
NAND2XL inst_cellmath__64_0_I515 (.Y(N1742), .A(N1627), .B(N1629));
NOR2XL inst_cellmath__64_0_I516 (.Y(N1743), .A(N1630), .B(N1632));
NAND2XL inst_cellmath__64_0_I517 (.Y(N1744), .A(N1630), .B(N1632));
NOR2XL inst_cellmath__64_0_I518 (.Y(N1745), .A(N1633), .B(N1635));
NAND2XL inst_cellmath__64_0_I519 (.Y(N1746), .A(N1633), .B(N1635));
NOR2XL inst_cellmath__64_0_I520 (.Y(N1747), .A(N1636), .B(N1638));
NAND2XL inst_cellmath__64_0_I521 (.Y(N1748), .A(N1636), .B(N1638));
NOR2XL inst_cellmath__64_0_I522 (.Y(N1749), .A(N1639), .B(N1641));
NAND2XL inst_cellmath__64_0_I523 (.Y(N1750), .A(N1639), .B(N1641));
NOR2XL inst_cellmath__64_0_I524 (.Y(N1751), .A(N1642), .B(N1644));
NAND2XL inst_cellmath__64_0_I525 (.Y(N1752), .A(N1642), .B(N1644));
NOR2XL inst_cellmath__64_0_I526 (.Y(N1753), .A(N1645), .B(N1647));
NAND2XL inst_cellmath__64_0_I527 (.Y(N1754), .A(N1645), .B(N1647));
NOR2XL inst_cellmath__64_0_I528 (.Y(N1755), .A(N1648), .B(N1650));
NAND2XL inst_cellmath__64_0_I529 (.Y(N1756), .A(N1648), .B(N1650));
AOI21XL inst_cellmath__64_0_I532 (.Y(N1759), .A0(N1730), .A1(N1728), .B0(N1729));
INVXL inst_cellmath__64_0_I1878 (.Y(N3721), .A(N1731));
INVXL inst_cellmath__64_0_I1879 (.Y(N3722), .A(N1732));
OAI21XL inst_cellmath__64_0_I540 (.Y(N1767), .A0(N3722), .A1(N1759), .B0(N3721));
AOI21XL inst_cellmath__64_0_I548 (.Y(N1775), .A0(N1734), .A1(N1767), .B0(N1733));
INVXL inst_cellmath__64_0_I1885 (.Y(N3728), .A(N1735));
INVXL inst_cellmath__64_0_I1886 (.Y(N3729), .A(N1736));
OAI21XL inst_cellmath__64_0_I560 (.Y(N1787), .A0(N3729), .A1(N1775), .B0(N3728));
AOI21XL inst_cellmath__64_0_I572 (.Y(N1799), .A0(N1738), .A1(N1787), .B0(N1737));
INVXL inst_cellmath__64_0_I1900 (.Y(N3743), .A(N1739));
INVXL inst_cellmath__64_0_I1901 (.Y(N3744), .A(N1740));
OAI21XL inst_cellmath__64_0_I588 (.Y(N1815), .A0(N3744), .A1(N1799), .B0(N3743));
AOI21XL inst_cellmath__64_0_I604 (.Y(N1831), .A0(N1742), .A1(N1815), .B0(N1741));
INVXL inst_cellmath__64_0_I1919 (.Y(N3762), .A(N1743));
INVXL inst_cellmath__64_0_I1920 (.Y(N3763), .A(N1744));
OAI21XL inst_cellmath__64_0_I624 (.Y(N1851), .A0(N3763), .A1(N1831), .B0(N3762));
AOI21XL inst_cellmath__64_0_I644 (.Y(N1871), .A0(N1746), .A1(N1851), .B0(N1745));
INVXL inst_cellmath__64_0_I1942 (.Y(N3785), .A(N1747));
INVXL inst_cellmath__64_0_I1943 (.Y(N3786), .A(N1748));
OAI21XL inst_cellmath__64_0_I668 (.Y(N1895), .A0(N3786), .A1(N1871), .B0(N3785));
AOI21XL inst_cellmath__64_0_I692 (.Y(N1919), .A0(N1750), .A1(N1895), .B0(N1749));
INVXL inst_cellmath__64_0_I1969 (.Y(N3812), .A(N1751));
INVXL inst_cellmath__64_0_I1970 (.Y(N3813), .A(N1752));
OAI21XL inst_cellmath__64_0_I720 (.Y(N1947), .A0(N3813), .A1(N1919), .B0(N3812));
AOI21XL inst_cellmath__64_0_I748 (.Y(N1975), .A0(N1754), .A1(N1947), .B0(N1753));
INVXL inst_cellmath__64_0_I2000 (.Y(N3843), .A(N1755));
INVXL inst_cellmath__64_0_I2001 (.Y(N3844), .A(N1756));
OAI21XL inst_cellmath__64_0_I780 (.Y(N2070), .A0(N3844), .A1(N1975), .B0(N3843));
NAND2BXL inst_cellmath__64_0_I787 (.Y(N2014), .AN(N1729), .B(N1730));
NAND2BXL inst_cellmath__64_0_I790 (.Y(N2017), .AN(N1731), .B(N1732));
NAND2BXL inst_cellmath__64_0_I793 (.Y(N2020), .AN(N1733), .B(N1734));
NAND2BXL inst_cellmath__64_0_I796 (.Y(N2023), .AN(N1735), .B(N1736));
NAND2BXL inst_cellmath__64_0_I799 (.Y(N2026), .AN(N1737), .B(N1738));
NAND2BXL inst_cellmath__64_0_I802 (.Y(N2029), .AN(N1739), .B(N1740));
NAND2BXL inst_cellmath__64_0_I805 (.Y(N2032), .AN(N1741), .B(N1742));
NAND2BXL inst_cellmath__64_0_I808 (.Y(N2035), .AN(N1743), .B(N1744));
NAND2BXL inst_cellmath__64_0_I811 (.Y(N2038), .AN(N1745), .B(N1746));
NAND2BXL inst_cellmath__64_0_I814 (.Y(N2041), .AN(N1747), .B(N1748));
NAND2BXL inst_cellmath__64_0_I817 (.Y(N2044), .AN(N1749), .B(N1750));
NAND2BXL inst_cellmath__64_0_I820 (.Y(N2047), .AN(N1751), .B(N1752));
NAND2BXL inst_cellmath__64_0_I823 (.Y(N2050), .AN(N1753), .B(N1754));
NAND2BXL inst_cellmath__64_0_I826 (.Y(N2053), .AN(N1755), .B(N1756));
XOR2XL inst_cellmath__64_0_I2976 (.Y(inst_cellmath__64_0_out0[0]), .A(N1609), .B(inst_cellmath__64_0_in2[0]));
XOR2XL inst_cellmath__64_0_I2353 (.Y(inst_cellmath__64_0_out0[1]), .A(N1728), .B(N2014));
XNOR2X1 inst_cellmath__64_0_I829 (.Y(inst_cellmath__64_0_out0[2]), .A(N1759), .B(N2017));
XOR2XL inst_cellmath__64_0_I2354 (.Y(inst_cellmath__64_0_out0[3]), .A(N1767), .B(N2020));
XNOR2X1 inst_cellmath__64_0_I831 (.Y(inst_cellmath__64_0_out0[4]), .A(N1775), .B(N2023));
XOR2XL inst_cellmath__64_0_I2355 (.Y(inst_cellmath__64_0_out0[5]), .A(N1787), .B(N2026));
XNOR2X1 inst_cellmath__64_0_I833 (.Y(inst_cellmath__64_0_out0[6]), .A(N1799), .B(N2029));
XOR2XL inst_cellmath__64_0_I2356 (.Y(inst_cellmath__64_0_out0[7]), .A(N1815), .B(N2032));
XNOR2X1 inst_cellmath__64_0_I835 (.Y(inst_cellmath__64_0_out0[8]), .A(N1831), .B(N2035));
XOR2XL inst_cellmath__64_0_I2357 (.Y(inst_cellmath__64_0_out0[9]), .A(N1851), .B(N2038));
XNOR2X1 inst_cellmath__64_0_I837 (.Y(inst_cellmath__64_0_out0[10]), .A(N1871), .B(N2041));
XOR2XL inst_cellmath__64_0_I2358 (.Y(inst_cellmath__64_0_out0[11]), .A(N1895), .B(N2044));
XNOR2X1 inst_cellmath__64_0_I839 (.Y(inst_cellmath__64_0_out0[12]), .A(N1919), .B(N2047));
XOR2XL inst_cellmath__64_0_I2977 (.Y(inst_cellmath__64_0_out0[13]), .A(N1947), .B(N2050));
XNOR2X1 inst_cellmath__64_0_I841 (.Y(inst_cellmath__64_0_out0[14]), .A(N1975), .B(N2053));
NOR2XL inst_cellmath__64_0_I844 (.Y(N2072), .A(N1651), .B(N1653));
XOR2XL inst_cellmath__64_0_I845 (.Y(N2073), .A(N1651), .B(N1653));
XNOR2X1 inst_cellmath__64_0_I847 (.Y(N2075), .A(N1654), .B(N1656));
XOR2XL inst_cellmath__64_0_I849 (.Y(N2077), .A(N1657), .B(N1659));
XNOR2X1 inst_cellmath__64_0_I851 (.Y(N2079), .A(N1660), .B(N1662));
XOR2XL inst_cellmath__64_0_I853 (.Y(N2081), .A(N1663), .B(N1665));
XNOR2X1 inst_cellmath__64_0_I855 (.Y(N2083), .A(N1666), .B(N1668));
XOR2XL inst_cellmath__64_0_I857 (.Y(N2085), .A(N1669), .B(N1671));
XNOR2X1 inst_cellmath__64_0_I859 (.Y(N2087), .A(N1672), .B(N1674));
XOR2XL inst_cellmath__64_0_I861 (.Y(N2089), .A(N1675), .B(N1677));
XNOR2X1 inst_cellmath__64_0_I863 (.Y(N2091), .A(N1678), .B(N1680));
XOR2XL inst_cellmath__64_0_I865 (.Y(N2093), .A(N1683), .B(N1681));
XNOR2X1 inst_cellmath__64_0_I867 (.Y(N2095), .A(N1684), .B(N1686));
XOR2XL inst_cellmath__64_0_I869 (.Y(N2097), .A(N1687), .B(N1689));
XNOR2X1 inst_cellmath__64_0_I871 (.Y(N2099), .A(N1690), .B(N1692));
XOR2XL inst_cellmath__64_0_I873 (.Y(N2101), .A(N1693), .B(N1695));
XNOR2X1 inst_cellmath__64_0_I875 (.Y(N2103), .A(N1698), .B(N1696));
XOR2XL inst_cellmath__64_0_I877 (.Y(N2105), .A(N1701), .B(N1699));
XNOR2X1 inst_cellmath__64_0_I879 (.Y(N2107), .A(N1704), .B(N1702));
XOR2XL inst_cellmath__64_0_I881 (.Y(N2109), .A(N1707), .B(N1705));
XNOR2X1 inst_cellmath__64_0_I883 (.Y(N2111), .A(N1710), .B(N1708));
XOR2XL inst_cellmath__64_0_I885 (.Y(N2113), .A(N1713), .B(N1711));
XNOR2X1 inst_cellmath__64_0_I887 (.Y(N2115), .A(N1714), .B(N1716));
XOR2XL inst_cellmath__64_0_I889 (.Y(N2117), .A(N1717), .B(N1719));
XNOR2X1 inst_cellmath__64_0_I891 (.Y(N2119), .A(N1720), .B(N1722));
XNOR2X1 inst_cellmath__64_0_I893 (.Y(N2121), .A(N1723), .B(N1725));
AOI21XL inst_cellmath__64_0_I896 (.Y(N2124), .A0(N2073), .A1(N2070), .B0(N2072));
OAI22XL inst_cellmath__64_0_I2361 (.Y(N2132), .A0(N2075), .A1(N2124), .B0(N1654), .B1(N1656));
AOI2BB2X1 inst_cellmath__64_0_I1859 (.Y(N2140), .A0N(N1657), .A1N(N1659), .B0(N2132), .B1(N2077));
OAI22XL inst_cellmath__64_0_I2363 (.Y(N2152), .A0(N2079), .A1(N2140), .B0(N1660), .B1(N1662));
AOI2BB2X1 inst_cellmath__64_0_I1860 (.Y(N2164), .A0N(N1663), .A1N(N1665), .B0(N2152), .B1(N2081));
OAI22XL inst_cellmath__64_0_I2365 (.Y(N2180), .A0(N2083), .A1(N2164), .B0(N1666), .B1(N1668));
AOI2BB2X1 inst_cellmath__64_0_I1861 (.Y(N2196), .A0N(N1669), .A1N(N1671), .B0(N2180), .B1(N2085));
OAI22XL inst_cellmath__64_0_I2367 (.Y(N2216), .A0(N2087), .A1(N2196), .B0(N1672), .B1(N1674));
AOI2BB2X1 inst_cellmath__64_0_I1862 (.Y(N2236), .A0N(N1675), .A1N(N1677), .B0(N2216), .B1(N2089));
OAI22XL inst_cellmath__64_0_I2369 (.Y(N2260), .A0(N2091), .A1(N2236), .B0(N1678), .B1(N1680));
AOI2BB2X1 inst_cellmath__64_0_I1863 (.Y(N2284), .A0N(N1683), .A1N(N1681), .B0(N2260), .B1(N2093));
OAI22XL inst_cellmath__64_0_I2371 (.Y(N2312), .A0(N2095), .A1(N2284), .B0(N1684), .B1(N1686));
AOI2BB2X1 inst_cellmath__64_0_I1864 (.Y(N2340), .A0N(N1687), .A1N(N1689), .B0(N2312), .B1(N2097));
OAI22XL inst_cellmath__64_0_I2373 (.Y(N2372), .A0(N2099), .A1(N2340), .B0(N1690), .B1(N1692));
AOI2BB2X1 inst_cellmath__64_0_I1865 (.Y(N2404), .A0N(N1693), .A1N(N1695), .B0(N2372), .B1(N2101));
OAI22XL inst_cellmath__64_0_I2375 (.Y(N2440), .A0(N2103), .A1(N2404), .B0(N1698), .B1(N1696));
AOI2BB2X1 inst_cellmath__64_0_I1866 (.Y(N2476), .A0N(N1701), .A1N(N1699), .B0(N2440), .B1(N2105));
OAI22XL inst_cellmath__64_0_I2377 (.Y(N2516), .A0(N2107), .A1(N2476), .B0(N1704), .B1(N1702));
AOI2BB2X1 inst_cellmath__64_0_I1867 (.Y(N2556), .A0N(N1707), .A1N(N1705), .B0(N2516), .B1(N2109));
OAI22XL inst_cellmath__64_0_I2379 (.Y(N2600), .A0(N2111), .A1(N2556), .B0(N1710), .B1(N1708));
AOI2BB2X1 inst_cellmath__64_0_I2380 (.Y(N2644), .A0N(N1713), .A1N(N1711), .B0(N2600), .B1(N2113));
OAI22XL inst_cellmath__64_0_I2382 (.Y(N2692), .A0(N2115), .A1(N2644), .B0(N1714), .B1(N1716));
AOI2BB2X1 inst_cellmath__64_0_I2383 (.Y(N2740), .A0N(N1717), .A1N(N1719), .B0(N2692), .B1(N2117));
OA22X1 inst_cellmath__64_0_I2386 (.Y(N4195), .A0(N2119), .A1(N2740), .B0(N1720), .B1(N1722));
XNOR2X1 inst_cellmath__64_0_I2387 (.Y(inst_cellmath__64_0_out0[15]), .A(N2070), .B(N2073));
XNOR2X1 inst_cellmath__64_0_I1649 (.Y(inst_cellmath__64_0_out0[16]), .A(N2124), .B(N2075));
XNOR2X1 inst_cellmath__64_0_I1650 (.Y(inst_cellmath__64_0_out0[17]), .A(N2132), .B(N2077));
XNOR2X1 inst_cellmath__64_0_I1651 (.Y(inst_cellmath__64_0_out0[18]), .A(N2140), .B(N2079));
XNOR2X1 inst_cellmath__64_0_I1652 (.Y(inst_cellmath__64_0_out0[19]), .A(N2152), .B(N2081));
XNOR2X1 inst_cellmath__64_0_I1653 (.Y(inst_cellmath__64_0_out0[20]), .A(N2164), .B(N2083));
XNOR2X1 inst_cellmath__64_0_I1654 (.Y(inst_cellmath__64_0_out0[21]), .A(N2180), .B(N2085));
XNOR2X1 inst_cellmath__64_0_I1655 (.Y(inst_cellmath__64_0_out0[22]), .A(N2196), .B(N2087));
XNOR2X1 inst_cellmath__64_0_I1656 (.Y(inst_cellmath__64_0_out0[23]), .A(N2216), .B(N2089));
XNOR2X1 inst_cellmath__64_0_I1657 (.Y(inst_cellmath__64_0_out0[24]), .A(N2236), .B(N2091));
XNOR2X1 inst_cellmath__64_0_I1658 (.Y(inst_cellmath__64_0_out0[25]), .A(N2260), .B(N2093));
XNOR2X1 inst_cellmath__64_0_I1659 (.Y(inst_cellmath__64_0_out0[26]), .A(N2284), .B(N2095));
XNOR2X1 inst_cellmath__64_0_I1660 (.Y(inst_cellmath__64_0_out0[27]), .A(N2312), .B(N2097));
XNOR2X1 inst_cellmath__64_0_I1661 (.Y(inst_cellmath__64_0_out0[28]), .A(N2340), .B(N2099));
XNOR2X1 inst_cellmath__64_0_I1662 (.Y(inst_cellmath__64_0_out0[29]), .A(N2372), .B(N2101));
XNOR2X1 inst_cellmath__64_0_I1663 (.Y(inst_cellmath__64_0_out0[30]), .A(N2404), .B(N2103));
XNOR2X1 inst_cellmath__64_0_I1664 (.Y(inst_cellmath__64_0_out0[31]), .A(N2440), .B(N2105));
XNOR2X1 inst_cellmath__64_0_I1665 (.Y(inst_cellmath__64_0_out0[32]), .A(N2476), .B(N2107));
XNOR2X1 inst_cellmath__64_0_I1666 (.Y(inst_cellmath__64_0_out0[33]), .A(N2516), .B(N2109));
XNOR2X1 inst_cellmath__64_0_I1667 (.Y(inst_cellmath__64_0_out0[34]), .A(N2556), .B(N2111));
XNOR2X1 inst_cellmath__64_0_I1668 (.Y(inst_cellmath__64_0_out0[35]), .A(N2600), .B(N2113));
XNOR2X1 inst_cellmath__64_0_I1669 (.Y(inst_cellmath__64_0_out0[36]), .A(N2644), .B(N2115));
XNOR2X1 inst_cellmath__64_0_I1670 (.Y(inst_cellmath__64_0_out0[37]), .A(N2692), .B(N2117));
XNOR2X1 inst_cellmath__64_0_I1671 (.Y(inst_cellmath__64_0_out0[38]), .A(N2740), .B(N2119));
XNOR2X1 inst_cellmath__64_0_I1672 (.Y(inst_cellmath__64_0_out0[39]), .A(N4195), .B(N2121));
endmodule

module cynw_cm_float_rcp_inst_cellmath__68_0_bdw1412651405_bdw (
	inst_cellmath__68_0_out0,
	inst_cellmath__68_0_in0,
	inst_cellmath__68_0_in1,
	inst_cellmath__68_0_in2
	); /* architecture "gate_level" */ 
output [22:0] inst_cellmath__68_0_out0;
input  inst_cellmath__68_0_in0;
input [39:17] inst_cellmath__68_0_in1;
input  inst_cellmath__68_0_in2;
MX2XL inst_cellmath__68_0_I46 (.Y(inst_cellmath__68_0_out0[0]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[17]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I47 (.Y(inst_cellmath__68_0_out0[1]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[18]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I48 (.Y(inst_cellmath__68_0_out0[2]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[19]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I49 (.Y(inst_cellmath__68_0_out0[3]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[20]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I50 (.Y(inst_cellmath__68_0_out0[4]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[21]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I51 (.Y(inst_cellmath__68_0_out0[5]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[22]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I52 (.Y(inst_cellmath__68_0_out0[6]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[23]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I53 (.Y(inst_cellmath__68_0_out0[7]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[24]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I54 (.Y(inst_cellmath__68_0_out0[8]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[25]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I55 (.Y(inst_cellmath__68_0_out0[9]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[26]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I56 (.Y(inst_cellmath__68_0_out0[10]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[27]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I57 (.Y(inst_cellmath__68_0_out0[11]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[28]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I58 (.Y(inst_cellmath__68_0_out0[12]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[29]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I59 (.Y(inst_cellmath__68_0_out0[13]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[30]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I60 (.Y(inst_cellmath__68_0_out0[14]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[31]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I61 (.Y(inst_cellmath__68_0_out0[15]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[32]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I62 (.Y(inst_cellmath__68_0_out0[16]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[33]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I63 (.Y(inst_cellmath__68_0_out0[17]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[34]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I64 (.Y(inst_cellmath__68_0_out0[18]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[35]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I65 (.Y(inst_cellmath__68_0_out0[19]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[36]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I66 (.Y(inst_cellmath__68_0_out0[20]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[37]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I67 (.Y(inst_cellmath__68_0_out0[21]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[38]), .S0(inst_cellmath__68_0_in0));
MX2XL inst_cellmath__68_0_I68 (.Y(inst_cellmath__68_0_out0[22]), .A(inst_cellmath__68_0_in2), .B(inst_cellmath__68_0_in1[39]), .S0(inst_cellmath__68_0_in0));
endmodule

/* CADENCE  uLTzSwjeohk= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



