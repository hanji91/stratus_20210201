/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 12:10:30 KST (+0900), Tuesday 29 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module float_div_cynw_cm_float_rcp_E8_M23_0_0 (
	a_sign,
	a_exp,
	a_man,
	x
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
output [36:0] x;
wire  inst_cellmath__9,
	inst_cellmath__17;
wire [8:0] inst_cellmath__19;
wire [7:0] inst_cellmath__20;
wire [8:0] inst_cellmath__22;
wire  inst_cellmath__29,
	inst_cellmath__30,
	inst_cellmath__33,
	inst_cellmath__34,
	inst_cellmath__38,
	inst_cellmath__42;
wire [15:0] inst_cellmath__48;
wire [18:0] inst_cellmath__51;
wire [24:0] inst_cellmath__60;
wire [39:0] inst_cellmath__62__W0, inst_cellmath__62__W1,
	inst_cellmath__63__W0, inst_cellmath__63__W1;
wire [39:0] inst_cellmath__64;
wire  inst_cellmath__67;
wire N447,N449,N450,N451,N452,N454,N456 
	,N477,N478,N479,N480,N481,N482,N483,N484 
	,N485,N486,N487,N488,N489,N490,N491,N492 
	,N493,N494,N495,N496,N497,N498,N499,N500 
	,N501,N3125,N3127,N3142,N3148,N3158,N3161,N3163 
	,N3167,N3169,N3173,N3179,N3183,N3209,N3233,N3237 
	,N3240,N3241,N3244,N3246,N3247,N3248,N3250,N3254 
	,N3256,N3289,N3292,N3295,N3320,N3326,N3328,N3330 
	,N3335,N3338,N3392,N3394,N3395,N3397,N3399,N3400 
	,N3402,N3403,N3404,N3410,N3411,N3412,N3413,N3414 
	,N3416,N3417,N3418,N3419,N3421,N3422,N3424,N3425 
	,N3426,N3427,N3428,N3429,N3430,N3432,N3433,N3434 
	,N3437,N3438,N3439,N3441,N3442,N3444,N3446,N3450 
	,N3451,N3452,N3453,N3454,N3455,N3456,N3457,N3458 
	,N3459,N3460,N3461,N3462,N3463,N3464,N3466,N3467 
	,N3468,N3470,N3471,N3473,N3474,N3475,N3478,N3480 
	,N3482,N3483,N3485,N3486,N3487,N3488,N3489,N3491 
	,N3494,N3496,N3498,N3499,N3500,N3501,N3502,N3503 
	,N3504,N3506,N3507,N3508,N3509,N3510,N3511,N3512 
	,N3517,N3518,N3521,N3523,N3525,N3526,N3528,N3529 
	,N3530,N3532,N3534,N3535,N3537,N3538,N3540,N3541 
	,N3542,N3544,N3545,N3546,N3547,N3548,N3549,N3550 
	,N3553,N3554,N3555,N3556,N3558,N3559,N3560,N3562 
	,N3564,N3565,N3568,N3569,N3570,N3571,N3574,N3575 
	,N3577,N3579,N3580,N3581,N3582,N3583,N3584,N3588 
	,N3589,N3590,N3591,N3592,N3593,N3594,N3596,N3597 
	,N3598,N3600,N3601,N3603,N3604,N3605,N3608,N3609 
	,N3611,N3612,N3615,N3617,N3618,N3619,N3620,N3621 
	,N3623,N3624,N3625,N3626,N3627,N3628,N3629,N3630 
	,N3631,N3632,N3633,N3634,N3637,N3638,N3640,N3641 
	,N3642,N3643,N3644,N3646,N3647,N3648,N3649,N3656 
	,N3657,N3659,N3661,N3662,N3663,N3664,N3666,N3668 
	,N3669,N3670,N3672,N3673,N3674,N3675,N3676,N3678 
	,N3679,N3680,N3681,N3682,N3683,N3684,N3685,N3686 
	,N3687,N3690,N3691,N3692,N3694,N3695,N3696,N3698 
	,N3699,N3700,N3702,N3703,N3704,N3705,N3706,N3708 
	,N3709,N3710,N3712,N3713,N3714,N3715,N3716,N3717 
	,N3718,N3719,N3720,N3722,N3723,N3724,N3725,N3726 
	,N3729,N3730,N3731,N3734,N3735,N3737,N3739,N3741 
	,N3742,N3743,N3744,N3747,N3749,N3750,N3751,N3753 
	,N3754,N3756,N3758,N3759,N3760,N3761,N3762,N3763 
	,N3765,N3766,N3767,N3768,N3771,N3772,N3774,N3775 
	,N4147,N4148,N4149,N4150,N4151,N4152,N4153,N4154 
	,N4155,N4156,N4157,N4158,N4161,N4162,N4163,N4164 
	,N4165,N4166,N4167,N4168,N4170,N4171,N4172,N4173 
	,N4175,N4176,N4177,N4178,N4179,N4180,N4181,N4182 
	,N4183,N4185,N4186,N4187,N4188,N4189,N4190,N4191 
	,N4192,N4193,N4194,N4196,N4198,N4199,N4201,N4202 
	,N4203,N4204,N4205,N4206,N4207,N4208,N4209,N4210 
	,N4212,N4213,N4215,N4216,N4217,N4218,N4220,N4221 
	,N4222,N4223,N4224,N4225,N4226,N4227,N4228,N4229 
	,N4230,N4231,N4232,N4234,N4235,N4237,N4238,N4239 
	,N4240,N4241,N4242,N4243,N4244,N4245,N4246,N4247 
	,N4249,N4250,N4251,N4252,N4254,N4255,N4256,N4257 
	,N4258,N4259,N4260,N4261,N4262,N4263,N4264,N4265 
	,N4266,N4267,N4268,N4269,N4270,N4271,N4272,N4274 
	,N4275,N4276,N4277,N4278,N4279,N4280,N4281,N4282 
	,N4284,N4285,N4286,N4287,N4288,N4290,N4291,N4292 
	,N4293,N4295,N4296,N4297,N4298,N4299,N4300,N4301 
	,N4303,N4304,N4305,N4306,N4307,N4308,N4310,N4311 
	,N4312,N4313,N4314,N4315,N4316,N4317,N4318,N4319 
	,N4320,N4321,N4322,N4323,N4325,N4326,N4327,N4328 
	,N4329,N4330,N4333,N4334,N4335,N4336,N4337,N4338 
	,N4339,N4340,N4341,N4344,N4346,N4347,N4348,N4349 
	,N4350,N4351,N4352,N4353,N4354,N4356,N4357,N4358 
	,N4360,N4361,N4362,N4363,N4364,N4365,N4366,N4367 
	,N4368,N4369,N4370,N4371,N4372,N4373,N4374,N4375 
	,N4376,N4377,N4379,N4380,N4381,N4382,N4383,N4385 
	,N4386,N4388,N4390,N4391,N4392,N4393,N4394,N4396 
	,N4397,N4398,N4399,N4400,N4401,N4402,N4403,N4404 
	,N4405,N4407,N4408,N4409,N4410,N4411,N4412,N4413 
	,N4414,N4415,N4416,N4418,N4419,N4420,N4421,N4422 
	,N4423,N4424,N4425,N4427,N4428,N4429,N4430,N4431 
	,N4433,N4434,N4435,N4436,N4437,N4438,N4439,N4440 
	,N4441,N4442,N4443,N4444,N4445,N4446,N4447,N4449 
	,N4450,N4451,N4452,N4453,N4454,N4455,N4456,N4457 
	,N4460,N4461,N4462,N4463,N4464,N4465,N4466,N4467 
	,N4468,N4469,N4470,N4471,N4472,N4473,N4476,N4477 
	,N4478,N4479,N4480,N4481,N4482,N4484,N4485,N4486 
	,N4487,N4489,N4490,N4491,N4492,N4494,N4495,N4496 
	,N4497,N4498,N4499,N4500,N4501,N4503,N4504,N4505 
	,N4506,N4507,N4508,N4509,N4510,N4512,N4513,N4515 
	,N4516,N4517,N4518,N4519,N4520,N4521,N4522,N4524 
	,N4525,N4526,N4527,N4528,N4529,N4530,N4531,N4532 
	,N4533,N4534,N4535,N4536,N4537,N4538,N4539,N4540 
	,N4541,N4542,N4543,N4544,N4546,N4547,N4548,N4549 
	,N4550,N4551,N4552,N4553,N4554,N4556,N4557,N4558 
	,N4559,N4560,N4561,N4563,N4564,N4565,N4566,N4568 
	,N4569,N4570,N4571,N4572,N4573,N4574,N4576,N4579 
	,N4580,N4581,N4582,N4583,N4584,N4585,N4586,N4588 
	,N4590,N4591,N4592,N4593,N4594,N4595,N4596,N4597 
	,N4598,N4599,N4600,N4601,N4602,N4603,N4605,N4606 
	,N4607,N4608,N4610,N4612,N4613,N4615,N4616,N4617 
	,N4618,N4619,N4621,N4622,N4623,N4624,N4626,N4627 
	,N4628,N4629,N4631,N4632,N4633,N4634,N4635,N4636 
	,N4637,N4638,N4639,N4640,N4641,N4642,N4643,N4644 
	,N4646,N4647,N4648,N4649,N4650,N4651,N4652,N4654 
	,N4656,N4657,N4659,N4660,N4661,N4662,N4663,N4664 
	,N4665,N4667,N4668,N4669,N4670,N4671,N4672,N4673 
	,N4674,N4675,N4676,N4677,N4678,N4680,N4681,N4682 
	,N4683,N4685,N4686,N4687,N4688,N4689,N4690,N4691 
	,N4692,N4694,N4695,N4696,N4697,N4698,N4700,N4701 
	,N4702,N4703,N4704,N4705,N4706,N4707,N4708,N4709 
	,N4711,N4712,N4713,N4714,N4715,N4716,N4717,N4718 
	,N4720,N4721,N4722,N4723,N4724,N4726,N4727,N4728 
	,N4729,N4732,N4733,N4734,N4735,N4736,N4738,N4739 
	,N4740,N4741,N4742,N4743,N4744,N4745,N4746,N4747 
	,N4749,N4750,N4752,N4753,N4754,N4755,N4756,N4758 
	,N4759,N4760,N4761,N4763,N4764,N4765,N4767,N4768 
	,N4770,N4771,N4772,N4773,N4774,N4776,N4777,N4778 
	,N4779,N4780,N4782,N4783,N4784,N4785,N4786,N4791 
	,N4792,N4793,N4794,N4796,N4797,N4798,N4799,N4800 
	,N4802,N4803,N4804,N4805,N4806,N4807,N4808,N4809 
	,N4810,N4812,N4813,N4814,N4815,N4816,N4817,N4818 
	,N4819,N4820,N4821,N4822,N4823,N4824,N4825,N4826 
	,N4828,N4829,N4830,N4831,N4833,N4834,N4835,N4836 
	,N4839,N4841,N4843,N4844,N4845,N4846,N4847,N4848 
	,N4849,N4850,N4851,N4852,N4854,N4855,N4856,N4857 
	,N4858,N4859,N4860,N4861,N4862,N4864,N4865,N4867 
	,N4868,N4869,N4871,N4872,N4873,N4875,N4876,N4877 
	,N4878,N4879,N4881,N4882,N4883,N4884,N4885,N4886 
	,N4887,N4888,N4889,N4890,N4891,N4892,N4894,N4895 
	,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4903 
	,N4905,N4906,N4907,N4908,N4909,N4910,N4911,N4912 
	,N4913,N4914,N4915,N4916,N4917,N4918,N4919,N4920 
	,N4922,N4923,N4924,N4925,N4926,N4927,N4928,N4929 
	,N4930,N4931,N4932,N4933,N4934,N4935,N4936,N4937 
	,N4938,N4939,N4941,N4942,N4944,N4945,N4947,N4948 
	,N4949,N4950,N4951,N4952,N4953,N4954,N4955,N4956 
	,N4957,N4958,N4961,N4962,N4963,N4964,N4965,N4966 
	,N4967,N4968,N4969,N4970,N4971,N4972,N4974,N4975 
	,N4977,N4978,N4979,N4980,N4981,N4982,N4983,N4984 
	,N4985,N4986,N4987,N4988,N4989,N4990,N4991,N4993 
	,N4994,N4995,N4996,N4997,N4998,N5000,N5001,N5002 
	,N5004,N5005,N5006,N5007,N5009,N5010,N5012,N5013 
	,N5014,N5015,N5016,N5017,N5018,N5019,N5020,N5021 
	,N5022,N5024,N5025,N5026,N5027,N5028,N5029,N5030 
	,N5031,N5032,N5035,N5036,N5037,N5039,N5040,N5041 
	,N5042,N5043,N5045,N5046,N5047,N5050,N5051,N5052 
	,N5053,N5054,N5055,N5056,N5057,N5058,N5059,N5060 
	,N5061,N5062,N5063,N5064,N5066,N5068,N5069,N5070 
	,N5071,N5072,N5073,N5074,N5075,N5076,N5077,N5078 
	,N5079,N5080,N5081,N5082,N5083,N5085,N5087,N5088 
	,N5089,N5090,N5091,N5093,N5094,N5095,N5096,N5097 
	,N5098,N5099,N5100,N5101,N5102,N5103,N5104,N5106 
	,N5107,N5108,N5109,N5110,N5111,N5112,N5113,N5115 
	,N5116,N5117,N5118,N5119,N5120,N5121,N5122,N5123 
	,N5124,N5125,N5126,N5127,N5128,N5129,N5131,N5132 
	,N5133,N5134,N5136,N5137,N5138,N5139,N5140,N5141 
	,N5142,N5143,N5145,N5146,N5147,N5148,N5149,N5150 
	,N5151,N5152,N5153,N5156,N5157,N5158,N5159,N5160 
	,N5161,N5163,N6174,N6176,N6178,N6179,N6181,N6182 
	,N6183,N6184,N6185,N6188,N6189,N6190,N6191,N6192 
	,N6195,N6196,N6197,N6198,N6199,N6200,N6201,N6202 
	,N6203,N6204,N6206,N6207,N6209,N6210,N6211,N6213 
	,N6214,N6216,N6217,N6218,N6220,N6222,N6223,N6224 
	,N6225,N6226,N6227,N6228,N6230,N6231,N6232,N6233 
	,N6234,N6235,N6237,N6238,N6239,N6241,N6242,N6243 
	,N6244,N6245,N6246,N6247,N6249,N6251,N6253,N6255 
	,N6256,N6257,N6258,N6259,N6260,N6262,N6264,N6265 
	,N6266,N6267,N6268,N6269,N6270,N6273,N6274,N6275 
	,N6276,N6277,N6278,N6279,N6281,N6283,N6284,N6285 
	,N6286,N6287,N6288,N6289,N6290,N6291,N6295,N6296 
	,N6297,N6298,N6299,N6301,N6302,N6304,N6305,N6306 
	,N6307,N6308,N6309,N6310,N6311,N6315,N6316,N6317 
	,N6318,N6319,N6320,N6321,N6323,N6324,N6326,N6327 
	,N6328,N6329,N6330,N6331,N6332,N6333,N6334,N6336 
	,N6337,N6339,N6341,N6342,N6344,N6345,N6347,N6348 
	,N6349,N6350,N6351,N6353,N6354,N6355,N6357,N6358 
	,N6359,N6360,N6361,N6362,N6363,N6365,N6367,N6369 
	,N6370,N6371,N6372,N6373,N6374,N6376,N6378,N6379 
	,N6380,N6381,N6382,N6383,N6385,N6386,N6387,N6389 
	,N6390,N6391,N6392,N6393,N6394,N6396,N6397,N6399 
	,N6401,N6402,N6403,N6404,N6405,N6407,N6408,N6409 
	,N6411,N6412,N6413,N6414,N6415,N6416,N6417,N6419 
	,N6420,N6421,N6422,N6423,N6424,N6425,N6427,N6428 
	,N6430,N6431,N6432,N6433,N6434,N6435,N6436,N6437 
	,N6438,N6440,N6442,N6444,N6445,N6446,N6447,N6449 
	,N6451,N6452,N6453,N6454,N6455,N6456,N6457,N6458 
	,N6459,N6464,N6465,N6466,N6467,N6468,N6469,N6470 
	,N6473,N6474,N6475,N6476,N6477,N6478,N6479,N6480 
	,N6482,N6483,N6484,N6486,N6488,N6489,N6490,N6491 
	,N6492,N6493,N6494,N6496,N6497,N6498,N6499,N6500 
	,N6501,N6502,N6503,N6505,N6507,N6508,N6509,N6510 
	,N6511,N6512,N6513,N6832,N6833,N6834,N6835,N6837 
	,N6839,N6840,N6841,N6842,N6843,N6844,N6845,N6846 
	,N6847,N6848,N6849,N6850,N6851,N6852,N6853,N6854 
	,N6855,N6856,N6857,N6859,N6860,N6861,N6863,N6864 
	,N6865,N6866,N6868,N6869,N6870,N6871,N6873,N6874 
	,N6875,N6876,N6877,N6878,N6880,N6881,N6882,N6883 
	,N6884,N6885,N6886,N6887,N6888,N6889,N6891,N6892 
	,N6893,N6894,N6895,N6896,N6897,N6899,N6900,N6901 
	,N6902,N6903,N6904,N6905,N6907,N6908,N6909,N6910 
	,N6911,N6912,N6913,N6914,N6916,N6917,N6918,N6919 
	,N6920,N6921,N6922,N6923,N6924,N6925,N6927,N6929 
	,N6931,N6932,N6933,N6934,N6935,N6936,N6937,N6939 
	,N6940,N6941,N6943,N6944,N6945,N6946,N6948,N6949 
	,N6950,N6951,N6952,N6953,N6954,N6955,N6956,N6957 
	,N6958,N6960,N6961,N6962,N6963,N6964,N6965,N6966 
	,N6968,N6969,N6970,N6971,N6972,N6974,N6975,N6976 
	,N6977,N6978,N6981,N6982,N6983,N6985,N6986,N6987 
	,N6988,N6989,N6990,N6992,N6994,N6995,N6996,N6997 
	,N6998,N6999,N7000,N7001,N7002,N7003,N7004,N7005 
	,N7006,N7007,N7009,N7010,N7011,N7012,N7013,N7014 
	,N7015,N7016,N7018,N7019,N7020,N7021,N7022,N7023 
	,N7025,N7026,N7028,N7029,N7031,N7032,N7034,N7035 
	,N7036,N7037,N7038,N7039,N7040,N7043,N7044,N7045 
	,N7046,N7047,N7048,N7049,N7050,N7051,N7052,N7054 
	,N7055,N7056,N7057,N7058,N7060,N7061,N7063,N7064 
	,N7065,N7066,N7067,N7068,N7069,N7071,N7072,N7073 
	,N7074,N7075,N7077,N7078,N7079,N7080,N7081,N7082 
	,N7083,N7084,N7085,N7086,N7087,N7088,N7089,N7090 
	,N7091,N7093,N7094,N7095,N7096,N7097,N7098,N7100 
	,N7101,N7102,N7103,N7104,N7105,N7106,N7107,N7108 
	,N7110,N7111,N7112,N7113,N7114,N7115,N7116,N7117 
	,N7118,N7120,N7121,N7122,N7123,N7125,N7127,N7128 
	,N7129,N7130,N7132,N7133,N7135,N7136,N7137,N7138 
	,N7140,N7141,N7142,N7143,N7145,N7146,N7147,N7148 
	,N7149,N7150,N7151,N7152,N7153,N7154,N7155,N7156 
	,N7157,N7158,N7159,N7160,N7161,N7162,N7164,N7165 
	,N7166,N7167,N7169,N7170,N7171,N7173,N7174,N7175 
	,N7176,N7178,N7179,N7180,N7181,N7182,N7183,N7184 
	,N7185,N7187,N7188,N7189,N7190,N7191,N7192,N7193 
	,N7194,N7196,N7197,N7198,N7199,N7200,N7202,N7203 
	,N7204,N7205,N7206,N7208,N7210,N7211,N7212,N7214 
	,N7215,N7216,N7217,N7219,N7220,N7221,N7222,N7223 
	,N7224,N7225,N7226,N7227,N7228,N7229,N7232,N7233 
	,N7234,N7235,N7236,N7237,N7238,N7240,N7241,N7243 
	,N7244,N7245,N7247,N7248,N7249,N7250,N7251,N7253 
	,N7254,N7255,N7256,N7257,N7258,N7259,N7260,N7261 
	,N7263,N7264,N7265,N7266,N7267,N7268,N7269,N7270 
	,N7271,N7272,N7274,N7275,N7276,N7277,N7279,N7281 
	,N7282,N7283,N7284,N7285,N7287,N7288,N7289,N7290 
	,N7291,N7292,N7293,N7294,N7295,N7296,N7298,N7299 
	,N7300,N7301,N7302,N7303,N7304,N7305,N7306,N7307 
	,N7308,N7309,N7310,N7311,N7312,N7313,N7315,N7316 
	,N7317,N7318,N7319,N7320,N7321,N7322,N7323,N7325 
	,N7326,N7327,N7328,N7330,N7331,N7333,N7334,N7335 
	,N7336,N7337,N7338,N7339,N7340,N7341,N7342,N7344 
	,N7345,N7346,N7347,N7348,N7349,N7350,N7351,N7352 
	,N7353,N7354,N7356,N7357,N7358,N7359,N7360,N7362 
	,N7363,N7365,N7366,N7367,N7368,N7369,N7370,N7371 
	,N7372,N7373,N7374,N7375,N7376,N7378,N7379,N7380 
	,N7381,N7382,N7383,N7384,N7385,N7386,N7387,N7388 
	,N7389,N7390,N7391,N7392,N7394,N7396,N7398,N7399 
	,N7401,N7402,N7404,N7405,N7406,N7407,N7408,N7409 
	,N7410,N7411,N7413,N7414,N7415,N7416,N7417,N7418 
	,N7419,N7420,N7421,N7422,N7423,N7424,N7427,N7428 
	,N7429,N7430,N7431,N7432,N7433,N7435,N7436,N7437 
	,N7439,N7440,N7441,N7442,N7444,N7445,N7446,N7449 
	,N7450,N7451,N7452,N7453,N7454,N7456,N7457,N7458 
	,N7459,N7460,N7463,N7464,N7465,N7466,N7467,N7468 
	,N7469,N7470,N7472,N7473,N7474,N7475,N7476,N7477 
	,N7479,N7480,N7481,N7483,N7484,N7485,N7486,N7487 
	,N7488,N7489,N7490,N7491,N7492,N7493,N7495,N7497 
	,N7498,N7499,N7500,N7501,N7502,N7503,N7504,N7505 
	,N7506,N7507,N7508,N7509,N7510,N7512,N7513,N7514 
	,N7515,N7516,N7517,N7518,N7519,N7520,N7522,N7523 
	,N7524,N7526,N7527,N7529,N7530,N7531,N7532,N7533 
	,N7534,N7535,N7536,N7538,N7539,N7540,N7541,N7542 
	,N7543,N7544,N7545,N7546,N7547,N7548,N7550,N7551 
	,N7553,N7554,N7555,N7556,N7558,N7559,N7560,N7561 
	,N7562,N7563,N7564,N7565,N7566,N7567,N7568,N7570 
	,N7571,N7572,N7573,N7574,N7575,N7576,N7577,N7578 
	,N7579,N7580,N7581,N7582,N7583,N7584,N7585,N7587 
	,N7588,N7589,N7590,N7591,N7593,N7594,N7595,N7596 
	,N7598,N7599,N7600,N7601,N7602,N7603,N7604,N7606 
	,N7607,N7608,N7609,N7610,N7611,N7612,N7613,N7614 
	,N7615,N7616,N7617,N7620,N7621,N7622,N7623,N7624 
	,N7625,N7626,N7627,N7629,N7630,N7631,N7632,N7633 
	,N7634,N7636,N7637,N7639,N7640,N7641,N7642,N7643 
	,N7644,N7645,N7646,N7647,N7648,N7650,N7651,N7652 
	,N7654,N7655,N7656,N7657,N7658,N7659,N7660,N7661 
	,N7662,N7663,N7664,N7665,N7666,N7667,N7668,N7669 
	,N7670,N7672,N7673,N7675,N7676,N7677,N7679,N7680 
	,N7681,N7682,N7683,N7684,N7685,N7686,N7689,N7690 
	,N7691,N7692,N7693,N7694,N7695,N7696,N7697,N7698 
	,N7699,N7700,N7702,N7703,N7705,N7706,N7707,N7708 
	,N7710,N7711,N7712,N8562,N8563,N8566,N8567,N8568 
	,N8570,N8572,N8574,N8575,N8576,N8578,N8579,N8581 
	,N8584,N8586,N8588,N8589,N8592,N8593,N8596,N8597 
	,N8598,N8600,N8601,N8602,N8604,N8605,N8606,N8607 
	,N8610,N8612,N8613,N8616,N8617,N8619,N8622,N8625 
	,N8630,N8631,N8632,N8634,N8635,N8636,N8638,N8639 
	,N8642,N8643,N8648,N8651,N8653,N8655,N8657,N8661 
	,N8662,N8664,N8665,N8667,N8668,N8670,N8671,N8674 
	,N8675,N8677,N8679,N8680,N8683,N8686,N8688,N8690 
	,N8691,N8695,N8696,N8698,N8705,N8707,N8708,N8711 
	,N8715,N8718,N8719,N8720,N8721,N8724,N8727,N8730 
	,N8731,N8733,N8734,N8736,N8738,N8741,N8743,N8745 
	,N8746,N8747,N8749,N8750,N8752,N8754,N8756,N8759 
	,N8760,N8762,N8764,N8767,N8768,N8769,N8770,N8771 
	,N8772,N8773,N8774,N8777,N8778,N8783,N8789,N8790 
	,N8792,N8793,N8795,N8796,N8797,N8802,N8803,N8805 
	,N8806,N8807,N8811,N8814,N8817,N8818,N8820,N8822 
	,N8823,N8824,N8826,N8828,N8830,N8831,N8833,N8835 
	,N8836,N8839,N8840,N8842,N8843,N8846,N8848,N8850 
	,N8854,N8857,N8859,N8861,N8862,N8863,N8866,N8867 
	,N8868,N8873,N8877,N8879,N8881,N8889,N8892,N8893 
	,N8894,N8897,N8898,N8901,N8903,N8909,N8911,N8913 
	,N8917,N8918,N8922,N8925,N8926,N8928,N8929,N8930 
	,N8931,N8933,N8934,N8939,N8940,N8942,N8944,N8946 
	,N8948,N8949,N8951,N8953,N8956,N8957,N8960,N8963 
	,N8964,N8967,N8969,N8970,N8971,N8976,N8978,N8980 
	,N8983,N8986,N8988,N8989,N8991,N8992,N8993,N8994 
	,N8998,N8999,N9003,N9004,N9006,N9007,N9008,N9009 
	,N9010,N9011,N9013,N9014,N9015,N9017,N9019,N9023 
	,N9024,N9026,N9029,N9030,N9032,N9034,N9035,N9038 
	,N9039,N9040,N9042,N9047,N9053,N9054,N9056,N9057 
	,N9059,N9060,N9061,N9064,N9065,N9068,N9070,N9071 
	,N9072,N9075,N9080,N9081,N9086,N9087,N9088,N9090 
	,N9092,N9094,N9096,N9098,N9100,N9103,N9108,N9110 
	,N9112,N9117,N9120,N9122,N9125,N9126,N9128,N9129 
	,N9130,N9133,N9140,N9142,N9147,N9150,N9154,N9156 
	,N9157,N9158,N9161,N9162,N9164,N9165,N9167,N9168 
	,N9170,N9172,N9174,N9176,N9179,N9180,N9182,N9183 
	,N9185,N9189,N9190,N9192,N9193,N9195,N9197,N9198 
	,N9199,N9202,N9203,N9206,N9207,N9209,N9210,N9211 
	,N9214,N9217,N9218,N9220,N9221,N9223,N9231,N9234 
	,N9235,N9236,N9237,N9239,N9240,N9242,N9244,N9246 
	,N9247,N9248,N9251,N9252,N9257,N9258,N9259,N9260 
	,N9262,N9263,N9265,N9267,N9268,N9273,N9282,N9283 
	,N9284,N9285,N9288,N9292,N9294,N9299,N9307,N9934 
	,N13558,N13732,N13738,N13744,N13745,N13748,N13752,N13754 
	,N13759,N13760,N13761,N13762,N13763,N13764,N13766,N13767 
	,N13772,N13782,N13786,N13788,N13789,N13791,N13795,N13797 
	,N13803,N13806,N13807,N13813,N13851,N26089,N26090,N26095 
	,N26096,N26097,N26100,N26104,N26108,N26111,N26140,N26143 
	,N26147,N26149,N26151,N26156,N26158,N26165,N26168,N26170 
	,N26198,N26200,N26203,N26206,N26211,N26213,N26214,N26216 
	,N26219,N26222,N26225,N26227,N26229,N26230,N26233,N26236 
	,N26240,N26243,N26246,N26247,N26250,N26253,N26260,N26263 
	,N26266,N26307,N26312,N26314,N26315,N26318,N26322,N26325 
	,N26327,N26330,N26333,N26335,N26338,N26340,N26341,N26344 
	,N26348,N26349,N26352,N26354,N26359,N26363,N26399,N26407 
	,N26412,N26415,N26417,N26419,N26436,N26439,N26444,N26449 
	,N26452,N26455,N26458,N26461,N26464,N26468,N26473,N26474 
	,N26479,N26481,N26483,N26486,N26489,N26490,N26493,N26496 
	,N26499,N26504,N26548,N26553,N26556,N26561,N26562,N26563 
	,N26565,N26579,N26581,N26583,N26585,N26587,N26590,N26593 
	,N26594,N26596,N26598,N26601,N26603,N26606,N26608,N26610 
	,N26611,N26615,N26616,N26619,N26621,N26624,N26626,N26627 
	,N26629,N26634,N26636,N26637,N26638,N26688,N26692,N26698 
	,N26703,N26710,N26737;
NAND2XL inst_cellmath__9_0_I235 (.Y(N3127), .A(a_exp[6]), .B(a_exp[5]));
AND4XL inst_cellmath__9_0_I16267 (.Y(N3125), .A(a_exp[4]), .B(a_exp[3]), .C(a_exp[2]), .D(a_exp[1]));
NAND3XL hyperpropagate_4_1_A_I6061 (.Y(N13813), .A(a_exp[7]), .B(a_exp[0]), .C(N3125));
NOR2XL hyperpropagate_4_1_A_I6062 (.Y(inst_cellmath__9), .A(N3127), .B(N13813));
NOR2XL inst_cellmath__15__5__I248 (.Y(N3148), .A(a_man[10]), .B(a_man[9]));
NOR2XL inst_cellmath__15__5__I249 (.Y(N3158), .A(a_man[8]), .B(a_man[7]));
NOR2XL inst_cellmath__15__5__I250 (.Y(N3169), .A(a_man[6]), .B(a_man[5]));
NOR2XL inst_cellmath__15__5__I251 (.Y(N3179), .A(a_man[4]), .B(a_man[3]));
INVX1 inst_cellmath__15__5__I252 (.Y(N3142), .A(a_man[2]));
OR4X1 inst_cellmath__15__5__I16268 (.Y(N3163), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4BX1 inst_cellmath__15__5__I16271 (.Y(N3167), .AN(N3142), .B(a_man[0]), .C(N3163), .D(a_man[1]));
OR4X1 inst_cellmath__15__5__I16269 (.Y(N3173), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 inst_cellmath__15__5__I16270 (.Y(N3183), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NAND4XL inst_cellmath__15__5__I5941 (.Y(N3161), .A(N3148), .B(N3169), .C(N3158), .D(N3179));
NOR4BX1 cynw_cm_float_rcp_I16272 (.Y(inst_cellmath__19[0]), .AN(N3167), .B(N3161), .C(N3173), .D(N3183));
INVXL cynw_cm_float_rcp_I16250 (.Y(N3209), .A(inst_cellmath__9));
NOR2XL cynw_cm_float_rcp_I16251 (.Y(inst_cellmath__29), .A(N3209), .B(inst_cellmath__19[0]));
NOR2BX1 cynw_cm_float_rcp_I5850 (.Y(x[31]), .AN(a_sign), .B(inst_cellmath__29));
INVXL cynw_cm_float_rcp_I5 (.Y(inst_cellmath__20[0]), .A(a_exp[0]));
INVXL cynw_cm_float_rcp_I6 (.Y(inst_cellmath__20[1]), .A(a_exp[1]));
INVXL cynw_cm_float_rcp_I7 (.Y(inst_cellmath__20[2]), .A(a_exp[2]));
INVXL cynw_cm_float_rcp_I8 (.Y(inst_cellmath__20[3]), .A(a_exp[3]));
INVXL cynw_cm_float_rcp_I9 (.Y(inst_cellmath__20[4]), .A(a_exp[4]));
INVXL cynw_cm_float_rcp_I10 (.Y(inst_cellmath__20[5]), .A(a_exp[5]));
INVXL cynw_cm_float_rcp_I11 (.Y(inst_cellmath__20[6]), .A(a_exp[6]));
INVXL cynw_cm_float_rcp_I12 (.Y(inst_cellmath__20[7]), .A(a_exp[7]));
AND2XL inst_cellmath__22_0_I269 (.Y(N3250), .A(inst_cellmath__20[0]), .B(inst_cellmath__19[0]));
NOR2XL inst_cellmath__22_0_I271 (.Y(N3246), .A(inst_cellmath__20[1]), .B(N3250));
NOR2XL inst_cellmath__22_0_I272 (.Y(N3256), .A(inst_cellmath__20[3]), .B(inst_cellmath__20[2]));
NAND2BXL inst_cellmath__22_0_I274 (.Y(N3240), .AN(inst_cellmath__20[2]), .B(N3246));
NAND2XL inst_cellmath__22_0_I275 (.Y(N3237), .A(N3256), .B(N3246));
NOR2XL inst_cellmath__22_0_I276 (.Y(N3247), .A(inst_cellmath__20[5]), .B(inst_cellmath__20[4]));
INVXL inst_cellmath__22_0_I277 (.Y(N3254), .A(inst_cellmath__20[6]));
NAND2XL inst_cellmath__22_0_I278 (.Y(N3233), .A(N3254), .B(N3247));
XOR2XL inst_cellmath__22_0_I282 (.Y(inst_cellmath__22[0]), .A(inst_cellmath__20[0]), .B(inst_cellmath__19[0]));
XNOR2X1 inst_cellmath__22_0_I5851 (.Y(inst_cellmath__22[1]), .A(N3250), .B(inst_cellmath__20[1]));
XOR2XL inst_cellmath__22_0_I285 (.Y(inst_cellmath__22[2]), .A(N3246), .B(inst_cellmath__20[2]));
XNOR2X1 inst_cellmath__22_0_I286 (.Y(inst_cellmath__22[3]), .A(N3240), .B(inst_cellmath__20[3]));
XNOR2X1 inst_cellmath__22_0_I5852 (.Y(inst_cellmath__22[4]), .A(N3237), .B(inst_cellmath__20[4]));
NOR2XL inst_cellmath__22_0_I289 (.Y(N3248), .A(inst_cellmath__20[4]), .B(N3237));
XOR2XL inst_cellmath__22_0_I290 (.Y(inst_cellmath__22[5]), .A(inst_cellmath__20[5]), .B(N3248));
XOR2XL inst_cellmath__22_0_I291 (.Y(N3241), .A(N3247), .B(N3254));
MXI2XL inst_cellmath__22_0_I292 (.Y(inst_cellmath__22[6]), .A(N3241), .B(N3254), .S0(N3237));
XNOR2X1 inst_cellmath__22_0_I293 (.Y(N3244), .A(N3233), .B(inst_cellmath__20[7]));
MX2XL inst_cellmath__22_0_I294 (.Y(inst_cellmath__22[7]), .A(N3244), .B(inst_cellmath__20[7]), .S0(N3237));
NOR4BX1 inst_cellmath__22_0_I5853 (.Y(inst_cellmath__22[8]), .AN(N3247), .B(inst_cellmath__20[6]), .C(N3237), .D(inst_cellmath__20[7]));
NOR3XL inst_cellmath__17__6__I297 (.Y(N3292), .A(inst_cellmath__22[2]), .B(inst_cellmath__22[3]), .C(inst_cellmath__22[5]));
NOR2XL inst_cellmath__17__6__I298 (.Y(N3295), .A(inst_cellmath__22[6]), .B(inst_cellmath__22[7]));
NOR4BX1 inst_cellmath__17__6__I5854 (.Y(N3289), .AN(N3295), .B(inst_cellmath__22[0]), .C(inst_cellmath__22[4]), .D(inst_cellmath__22[1]));
AO21XL cynw_cm_float_rcp_I5855 (.Y(inst_cellmath__17), .A0(N3292), .A1(N3289), .B0(inst_cellmath__22[8]));
NAND2XL cynw_cm_float_rcp_I303 (.Y(inst_cellmath__30), .A(N3209), .B(inst_cellmath__17));
OAI2BB1X1 cynw_cm_float_rcp_I5856 (.Y(N447), .A0N(inst_cellmath__9), .A1N(inst_cellmath__19[0]), .B0(inst_cellmath__30));
NOR2XL inst_cellmath__34_0_I307 (.Y(N3335), .A(a_exp[0]), .B(a_exp[1]));
NOR2XL inst_cellmath__34_0_I308 (.Y(N3338), .A(a_exp[7]), .B(a_exp[6]));
NOR2XL inst_cellmath__34_0_I309 (.Y(N3326), .A(a_exp[5]), .B(a_exp[4]));
NOR2XL inst_cellmath__34_0_I310 (.Y(N3330), .A(a_exp[3]), .B(a_exp[2]));
NAND4XL inst_cellmath__34_0_I311 (.Y(N3328), .A(N3335), .B(N3326), .C(N3338), .D(N3330));
NOR2XL cynw_cm_float_rcp_I16252 (.Y(inst_cellmath__34), .A(N3328), .B(inst_cellmath__29));
OR2XL inst_cellmath__42__9__I313 (.Y(inst_cellmath__38), .A(inst_cellmath__29), .B(inst_cellmath__34));
INVXL cynw_cm_float_rcp_I16253 (.Y(N3320), .A(inst_cellmath__29));
AND2XL cynw_cm_float_rcp_I16254 (.Y(inst_cellmath__33), .A(N3320), .B(N447));
NOR2XL inst_cellmath__42__9__I314 (.Y(inst_cellmath__42), .A(inst_cellmath__38), .B(inst_cellmath__33));
MX2XL inst_cellmath__43_0_I316 (.Y(x[23]), .A(inst_cellmath__38), .B(inst_cellmath__22[0]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I317 (.Y(x[24]), .A(inst_cellmath__38), .B(inst_cellmath__22[1]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I318 (.Y(x[25]), .A(inst_cellmath__38), .B(inst_cellmath__22[2]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I319 (.Y(x[26]), .A(inst_cellmath__38), .B(inst_cellmath__22[3]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I320 (.Y(x[27]), .A(inst_cellmath__38), .B(inst_cellmath__22[4]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I321 (.Y(x[28]), .A(inst_cellmath__38), .B(inst_cellmath__22[5]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I322 (.Y(x[29]), .A(inst_cellmath__38), .B(inst_cellmath__22[6]), .S0(inst_cellmath__42));
MX2XL inst_cellmath__43_0_I323 (.Y(x[30]), .A(inst_cellmath__38), .B(inst_cellmath__22[7]), .S0(inst_cellmath__42));
OR4X1 cynw_cm_float_rcp_I16255 (.Y(N26688), .A(inst_cellmath__29), .B(inst_cellmath__34), .C(inst_cellmath__19[0]), .D(inst_cellmath__33));
INVXL cynw_cm_float_rcp_I16256 (.Y(inst_cellmath__67), .A(N26688));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I16174 (.Y(N4911), .A(a_man[22]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I1166 (.Y(N4634), .A(a_man[21]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I920 (.Y(N4896), .A(a_man[20]));
CLKINVX8 inst_noninc_a_cellmath__55_2WWMM_I775 (.Y(N4533), .A(a_man[19]));
CLKINVX8 inst_noninc_a_cellmath__55_2WWMM_I651 (.Y(N4516), .A(a_man[17]));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I5794 (.Y(N13759), .A(N4516));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I5795 (.Y(N13760), .A(N13759));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I691 (.Y(N4350), .A(a_man[18]));
CLKINVX6 inst_noninc_a_cellmath__55_2WWMM_I694 (.Y(N5015), .A(N4350));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I695 (.Y(N4314), .A(N5015));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I5779 (.Y(N13744), .A(a_man[16]));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I656 (.Y(N4421), .A0(a_man[16]), .A1(N4516), .B0(N13744), .B1(a_man[17]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I657 (.Y(N4739), .A(N4421));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I658 (.Y(N4613), .A(N4739));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5796 (.Y(N13761), .A(N4613));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5801 (.Y(N13766), .A(N13761));
CLKINVX8 inst_noninc_a_cellmath__55_2WWMM_I5780 (.Y(N13745), .A(N13744));
NOR2X4 inst_noninc_a_cellmath__55_2WWMM_I16276 (.Y(N4479), .A(a_man[17]), .B(N13745));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5802 (.Y(N13767), .A(N5015));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5817 (.Y(N13782), .A(N13767));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1289 (.Y(N4576), .A0(N4314), .A1(N13766), .B0(N4479), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1494 (.Y(N4199), .A0(N4533), .A1(N13760), .B0(N4576), .B1(a_man[19]));
NAND2X6 inst_noninc_a_cellmath__55_2WWMM_I661 (.Y(N4869), .A(N13760), .B(N13744));
CLKINVX12 inst_noninc_a_cellmath__55_2WWMM_I5824 (.Y(N13789), .A(N4314));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5838 (.Y(N13803), .A(N13789));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I852 (.Y(N4276), .A0(N4869), .A1(N13782), .B0(N13803), .B1(N13760));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I707 (.Y(N4826), .A(N4350));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5841 (.Y(N13806), .A(N13789));
NOR2X4 inst_noninc_a_cellmath__55_2WWMM_I669 (.Y(N4736), .A(N13744), .B(N13760));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I833 (.Y(N4344), .A0(N13760), .A1(N4826), .B0(N13806), .B1(N4736));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I892 (.Y(N4651), .A0(N4533), .A1(N4276), .B0(N4344), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1542 (.Y(N4955), .A0(N4896), .A1(N4199), .B0(N4651), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1290 (.Y(N4225), .A0(N4314), .A1(N4869), .B0(N4736), .B1(N13782));
NAND2X4 inst_noninc_a_cellmath__55_2WWMM_I673 (.Y(N4166), .A(N13745), .B(a_man[17]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I5842 (.Y(N13807), .A(N13789));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5821 (.Y(N13786), .A(N13767));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1070 (.Y(N4706), .A0(N4166), .A1(N13807), .B0(a_man[17]), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1330 (.Y(N4626), .A0(N4533), .A1(N4225), .B0(N4706), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I732 (.Y(N4501), .A0(N13760), .A1(N4314), .B0(a_man[17]), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I6014 (.Y(N4271), .A0(N13760), .A1(N4314), .B0(N4736), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1268 (.Y(N4376), .A0(N4533), .A1(N4501), .B0(N4271), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1379 (.Y(N4581), .A0(N4896), .A1(N4626), .B0(N4376), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1594 (.Y(N4596), .A0(N4634), .A1(N4955), .B0(N4581), .B1(a_man[21]));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5826 (.Y(N13791), .A(N13789));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I5880 (.Y(N4619), .A(N13791), .B(N4166));
INVX3 inst_noninc_a_cellmath__55_2WWMM_I5830 (.Y(N13795), .A(N13789));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I740 (.Y(N5163), .A(N13795), .B(N4479));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5886 (.Y(N4816), .A0(N4533), .A1(N4619), .B0(N5163), .B1(a_man[19]));
NOR2X1 inst_noninc_a_cellmath__55_2WWMM_I731 (.Y(N4849), .A(N4826), .B(a_man[17]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I864 (.Y(N4413), .A(N13782), .B(N4869));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1041 (.Y(N4319), .A0(N4849), .A1(N4533), .B0(N4413), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5890 (.Y(N4993), .A0(N4896), .A1(N4816), .B0(N4319), .B1(a_man[20]));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5823 (.Y(N13788), .A(N13767));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I915 (.Y(N4852), .A0(N4533), .A1(N13788), .B0(N4849), .B1(a_man[19]));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I756 (.Y(N4644), .A(N13791), .B(N4479));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I817 (.Y(N4848), .A(N4533), .B(N4644));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I963 (.Y(N4808), .A0(N4896), .A1(N4852), .B0(N4848), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5893 (.Y(N4155), .A0(N4634), .A1(N4993), .B0(N4808), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5901 (.Y(N497), .A0(N4911), .A1(N4596), .B0(N4155), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2590 (.CO(N9133), .S(N8976), .A(1'B1), .B(N497));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I774 (.Y(N4252), .A0(N13803), .A1(N4479), .B0(N4869), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1495 (.Y(N4419), .A0(N4314), .A1(N4533), .B0(N4252), .B1(a_man[19]));
NAND2X1 inst_noninc_a_cellmath__55_2WWMM_I978 (.Y(N4341), .A(N13791), .B(N13760));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I819 (.Y(N5088), .A(N13803), .B(N13760));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1436 (.Y(N5029), .A0(N4533), .A1(N4341), .B0(N5088), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1543 (.Y(N4156), .A0(N4896), .A1(N4419), .B0(N5029), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5894 (.Y(N4847), .A0(N4533), .A1(N4314), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1269 (.Y(N4603), .A0(N4533), .A1(N4849), .B0(N4341), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5895 (.Y(N4803), .A0(N4896), .A1(N4847), .B0(N4603), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5899 (.Y(N4817), .A0(N4634), .A1(N4156), .B0(N4803), .B1(a_man[21]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I711 (.Y(N4349), .A(N4826), .B(N4736));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1114 (.Y(N5041), .A0(N4533), .A1(N4349), .B0(N5163), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1160 (.Y(N4198), .A0(N4896), .A1(N5041), .B0(a_man[19]), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I916 (.Y(N5074), .A(a_man[19]), .B(N13788));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I755 (.Y(N4968), .A(N4826), .B(N4869));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I818 (.Y(N4279), .A(N4533), .B(N4968));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I964 (.Y(N5030), .A0(N4896), .A1(N5074), .B0(N4279), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1215 (.Y(N4373), .A0(N4634), .A1(N4198), .B0(N5030), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5902 (.Y(N498), .A0(N4911), .A1(N4817), .B0(N4373), .B1(a_man[22]));
INVXL hap1_A_I16277 (.Y(N8771), .A(N498));
NOR2XL cynw_cm_float_rcp_I16257 (.Y(N9251), .A(N9133), .B(N8771));
NAND2XL cynw_cm_float_rcp_I16258 (.Y(N8670), .A(N9133), .B(N8771));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1555 (.Y(N4439), .A(a_man[20]), .B(N4279));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1556 (.Y(N4429), .A(N4439), .B(N4634));
OR2X1 inst_cellmath__62_0_I5915 (.Y(N6347), .A(a_man[22]), .B(N4429));
CLKINVX16 inst_cellmath__60_0_I332 (.Y(N3702), .A(a_man[9]));
CLKINVX6 inst_cellmath__60_0_I334 (.Y(N3432), .A(a_man[11]));
NOR2X1 inst_cellmath__60_0_I406 (.Y(N3418), .A(N3702), .B(N3432));
CLKINVX6 inst_cellmath__60_0_I339 (.Y(N3538), .A(a_man[14]));
CLKINVX6 inst_cellmath__60_0_I329 (.Y(N3412), .A(a_man[6]));
NOR2X1 inst_cellmath__60_0_I385 (.Y(N3414), .A(N3538), .B(N3412));
CLKINVX12 inst_cellmath__60_0_I16246 (.Y(N3611), .A(a_man[8]));
CLKINVX8 inst_cellmath__60_0_I336 (.Y(N3462), .A(a_man[12]));
NOR2XL inst_cellmath__60_0_I400 (.Y(N3716), .A(N3611), .B(N3462));
ADDFX1 inst_cellmath__60_0_I466 (.CO(N3558), .S(N3470), .A(N3418), .B(N3414), .CI(N3716));
CLKINVX12 inst_cellmath__60_0_I330 (.Y(N3446), .A(a_man[7]));
NOR2X1 inst_cellmath__60_0_I392 (.Y(N3672), .A(N3446), .B(N3462));
NOR2X1 inst_cellmath__60_0_I399 (.Y(N3544), .A(N3611), .B(N3432));
CLKINVX4 inst_cellmath__60_0_I16245 (.Y(N3456), .A(a_man[5]));
NOR2XL inst_cellmath__60_0_I375 (.Y(N3422), .A(N3456), .B(N3538));
ADDFXL inst_cellmath__60_0_I16138 (.CO(N3656), .S(N26349), .A(N3672), .B(N3544), .CI(N3422));
CLKINVX8 inst_cellmath__60_0_I333 (.Y(N3399), .A(a_man[10]));
NOR2XL inst_cellmath__60_0_I398 (.Y(N3759), .A(N3611), .B(N3399));
CLKINVX6 inst_cellmath__60_0_I338 (.Y(N3496), .A(a_man[13]));
NOR2XL inst_cellmath__60_0_I374 (.Y(N3638), .A(N3456), .B(N3496));
OR2XL inst_cellmath__60_0_I16132 (.Y(N26325), .A(N3759), .B(N3638));
CLKINVX6 inst_cellmath__60_0_I326 (.Y(N3503), .A(a_man[4]));
CLKINVX6 cynw_cm_float_rcp_I25 (.Y(inst_cellmath__48[15]), .A(a_man[15]));
CLKINVX4 inst_cellmath__60_0_I340 (.Y(N3571), .A(inst_cellmath__48[15]));
OR2XL inst_cellmath__60_0_I16125 (.Y(N26348), .A(N3503), .B(N3571));
NOR2X2 inst_cellmath__60_0_I383 (.Y(N3458), .A(N3462), .B(N3412));
NOR2X2 inst_cellmath__60_0_I391 (.Y(N3498), .A(N3446), .B(N3432));
NOR2X1 inst_cellmath__60_0_I364 (.Y(N3646), .A(N3503), .B(N3538));
ADDFXL inst_cellmath__60_0_I16133 (.CO(N26352), .S(N26338), .A(N3458), .B(N3498), .CI(N3646));
ADDFX1 inst_cellmath__60_0_I16139 (.CO(N3437), .S(N26315), .A(N26325), .B(N26348), .CI(N26352));
ADDFXL inst_cellmath__60_0_I468 (.CO(N3502), .S(N3425), .A(N3470), .B(N3656), .CI(N3437));
OR2XL inst_cellmath__60_0_I376 (.Y(N3601), .A(N3456), .B(N3571));
NOR2XL inst_cellmath__60_0_I393 (.Y(N3450), .A(N3446), .B(N3496));
NOR2X1 inst_cellmath__60_0_I405 (.Y(N3634), .A(N3702), .B(N3399));
INVXL inst_cellmath__60_0_I411 (.Y(N3556), .A(N3399));
NOR2XL inst_cellmath__60_0_I384 (.Y(N3630), .A(N3412), .B(N3496));
ADDFX1 inst_cellmath__60_0_I16137 (.CO(N3482), .S(N26322), .A(N3634), .B(N3556), .CI(N3630));
ADDFX1 inst_cellmath__60_0_I467 (.CO(N3725), .S(N3640), .A(N3601), .B(N3450), .CI(N3482));
NOR2X2 inst_cellmath__60_0_I412 (.Y(N3501), .A(N3399), .B(N3432));
INVX1 inst_cellmath__60_0_I417 (.Y(N3648), .A(N3432));
NOR2XL inst_cellmath__60_0_I394 (.Y(N3620), .A(N3446), .B(N3538));
ADDFX1 inst_cellmath__60_0_I470 (.CO(N3454), .S(N3758), .A(N3501), .B(N3648), .CI(N3620));
NOR2X1 inst_cellmath__60_0_I401 (.Y(N3487), .A(N3611), .B(N3496));
NOR2X1 inst_cellmath__60_0_I5771 (.Y(N13732), .A(N3702), .B(N3462));
OR2XL inst_cellmath__60_0_I386 (.Y(N3690), .A(N3412), .B(N3571));
ADDFXL inst_cellmath__60_0_I471 (.CO(N3626), .S(N3542), .A(N3487), .B(N13732), .CI(N3690));
ADDFHXL inst_cellmath__60_0_I472 (.CO(N3410), .S(N3715), .A(N3558), .B(N3758), .CI(N3542));
ADDFHX1 inst_cellmath__60_0_I473 (.CO(N3580), .S(N3486), .A(N3502), .B(N3725), .CI(N3715));
NOR2XL inst_cellmath__60_0_I408 (.Y(N3750), .A(N3702), .B(N3496));
NOR2XL inst_cellmath__60_0_I413 (.Y(N3676), .A(N3399), .B(N3462));
NOR2XL inst_cellmath__60_0_I402 (.Y(N3664), .A(N3611), .B(N3538));
ADDFX1 inst_cellmath__60_0_I474 (.CO(N3743), .S(N3663), .A(N3750), .B(N3676), .CI(N3664));
OR2XL inst_cellmath__60_0_I395 (.Y(N3774), .A(N3446), .B(N3571));
ADDFX1 inst_cellmath__60_0_I475 (.CO(N3529), .S(N3444), .A(N3454), .B(N3774), .CI(N3626));
ADDFX1 inst_cellmath__60_0_I476 (.CO(N3700), .S(N3609), .A(N3663), .B(N3410), .CI(N3444));
NOR2XL inst_cellmath__60_0_I540 (.Y(N3559), .A(N3580), .B(N3609));
NAND2X1 inst_cellmath__60_0_I541 (.Y(N3642), .A(N3580), .B(N3609));
NAND2BXL inst_cellmath__60_0_I600 (.Y(N3491), .AN(N3559), .B(N3642));
INVXL inst_cellmath__60_0_I404 (.Y(N3687), .A(N3702));
CLKINVX6 inst_cellmath__60_0_I341 (.Y(N3603), .A(a_man[3]));
NOR2X1 inst_cellmath__60_0_I353 (.Y(N3706), .A(N3603), .B(N3538));
ADDHX1 inst_cellmath__60_0_I16127 (.CO(N26340), .S(N26327), .A(N3687), .B(N3706));
OR2XL inst_cellmath__60_0_I16124 (.Y(N26335), .A(N3603), .B(N3571));
NOR2X4 inst_cellmath__60_0_I390 (.Y(N3722), .A(N3446), .B(N3399));
NOR2X4 inst_cellmath__60_0_I397 (.Y(N3591), .A(N3611), .B(N3702));
NOR2X2 inst_cellmath__60_0_I363 (.Y(N3473), .A(N3503), .B(N3496));
ADDFHXL inst_cellmath__60_0_I16128 (.CO(N26307), .S(N26354), .A(N3722), .B(N3591), .CI(N3473));
ADDFHXL inst_cellmath__60_0_I16134 (.CO(N26318), .S(N26363), .A(N26340), .B(N26335), .CI(N26307));
ADDFHXL inst_cellmath__60_0_I16140 (.CO(N3604), .S(N26341), .A(N26349), .B(N26322), .CI(N26318));
ADDFHXL inst_cellmath__60_0_I469 (.CO(N3678), .S(N3590), .A(N3604), .B(N3640), .CI(N3425));
NAND2X4 inst_cellmath__60_0_I539 (.Y(N3471), .A(N3678), .B(N3486));
XNOR2X1 inst_cellmath__60_0_I16131 (.Y(N26312), .A(N3759), .B(N3638));
NOR2XL inst_cellmath__60_0_I373 (.Y(N3468), .A(N3456), .B(N3462));
NOR2XL inst_cellmath__60_0_I382 (.Y(N3682), .A(N3412), .B(N3432));
NOR2XL inst_cellmath__60_0_I389 (.Y(N3553), .A(N3446), .B(N3702));
NOR2XL inst_cellmath__60_0_I352 (.Y(N3535), .A(N3603), .B(N3496));
ADDHX1 inst_cellmath__60_0_I446 (.CO(N3666), .S(N3581), .A(N3553), .B(N3535));
ADDFX1 inst_cellmath__60_0_I16129 (.CO(N26333), .S(N3433), .A(N3468), .B(N3682), .CI(N3666));
ADDFX1 inst_cellmath__60_0_I16135 (.CO(N26344), .S(N26330), .A(N26338), .B(N26312), .CI(N26333));
ADDFHXL inst_cellmath__60_0_I16141 (.CO(N3775), .S(N3694), .A(N26344), .B(N26315), .CI(N26341));
NAND2X2 inst_cellmath__60_0_I537 (.Y(N3695), .A(N3775), .B(N3590));
NAND2X4 inst_cellmath__60_0_I560 (.Y(N3463), .A(N3471), .B(N3695));
NOR2XL inst_cellmath__60_0_I362 (.Y(N3698), .A(N3503), .B(N3462));
NOR2XL inst_cellmath__60_0_I372 (.Y(N3691), .A(N3456), .B(N3432));
NOR2XL inst_cellmath__60_0_I381 (.Y(N3507), .A(N3412), .B(N3399));
ADDFX1 inst_cellmath__60_0_I16126 (.CO(N26314), .S(N3744), .A(N3698), .B(N3691), .CI(N3507));
ADDFXL inst_cellmath__60_0_I16130 (.CO(N26359), .S(N3598), .A(N26327), .B(N26354), .CI(N26314));
ADDFHXL inst_cellmath__60_0_I16136 (.CO(N3709), .S(N3619), .A(N26359), .B(N26363), .CI(N26330));
NAND2X4 inst_cellmath__60_0_I16142 (.Y(N3521), .A(N3709), .B(N3694));
INVXL inst_cellmath__60_0_I396 (.Y(N3641), .A(N3611));
NOR2XL inst_cellmath__60_0_I351 (.Y(N3749), .A(N3603), .B(N3462));
ADDHX1 inst_cellmath__60_0_I442 (.CO(N3761), .S(N3681), .A(N3641), .B(N3749));
NOR2XL inst_cellmath__60_0_I380 (.Y(N3729), .A(N3412), .B(N3702));
NOR2XL inst_cellmath__60_0_I388 (.Y(N3772), .A(N3446), .B(N3611));
NOR2XL inst_cellmath__60_0_I361 (.Y(N3525), .A(N3503), .B(N3432));
ADDFX1 inst_cellmath__60_0_I443 (.CO(N3547), .S(N3457), .A(N3729), .B(N3772), .CI(N3525));
ADDFX1 inst_cellmath__60_0_I448 (.CO(N3612), .S(N3532), .A(N3581), .B(N3761), .CI(N3547));
ADDFXL inst_cellmath__60_0_I454 (.CO(N3464), .S(N3771), .A(N3433), .B(N3612), .CI(N3598));
NAND2X2 inst_noninc_a_cellmath__55_2WWMM_I16168 (.Y(N3739), .A(N3464), .B(N3619));
NAND2X4 inst_cellmath__60_0_I558 (.Y(N3512), .A(N3739), .B(N3521));
NOR2X1 inst_cellmath__60_0_I577 (.Y(N3742), .A(N3463), .B(N3512));
NOR2XL inst_cellmath__60_0_I360 (.Y(N3741), .A(N3503), .B(N3399));
NOR2XL inst_cellmath__60_0_I370 (.Y(N3735), .A(N3456), .B(N3702));
INVXL inst_cellmath__60_0_I387 (.Y(N3434), .A(N3446));
NOR2XL inst_cellmath__60_0_I349 (.Y(N3416), .A(N3603), .B(N3399));
ADDHX1 inst_cellmath__60_0_I16219 (.CO(N26598), .S(N26583), .A(N3434), .B(N3416));
ADDFX1 inst_cellmath__60_0_I16223 (.CO(N3428), .S(N26626), .A(N3741), .B(N3735), .CI(N26598));
NOR2XL inst_cellmath__60_0_I379 (.Y(N3562), .A(N3412), .B(N3611));
NOR2XL inst_cellmath__60_0_I350 (.Y(N3583), .A(N3603), .B(N3432));
ADDHX1 inst_cellmath__60_0_I16222 (.CO(N3643), .S(N26601), .A(N3562), .B(N3583));
NOR2XL inst_cellmath__60_0_I371 (.Y(N3517), .A(N3456), .B(N3399));
ADDFX1 inst_cellmath__60_0_I444 (.CO(N3718), .S(N3628), .A(N3643), .B(N3517), .CI(N3681));
ADDFX1 inst_cellmath__60_0_I445 (.CO(N3489), .S(N3413), .A(N3428), .B(N3457), .CI(N3628));
ADDFX1 inst_cellmath__60_0_I449 (.CO(N3400), .S(N3703), .A(N3718), .B(N3744), .CI(N3532));
NAND2X1 inst_cellmath__60_0_I531 (.Y(N3574), .A(N3400), .B(N3771));
OAI2BB1X1 inst_cellmath__60_0_I5868 (.Y(N3565), .A0N(N3489), .A1N(N3703), .B0(N3574));
NOR2XL inst_cellmath__60_0_I16247 (.Y(N3568), .A(N3456), .B(N3611));
NOR2XL inst_cellmath__60_0_I378 (.Y(N3395), .A(N3412), .B(N3446));
NOR2XL inst_cellmath__60_0_I359 (.Y(N3577), .A(N3503), .B(N3702));
ADDFX1 inst_cellmath__60_0_I16220 (.CO(N26621), .S(N26608), .A(N3395), .B(N3568), .CI(N3577));
ADDFX1 inst_cellmath__60_0_I16224 (.CO(N3593), .S(N26596), .A(N26601), .B(N26621), .CI(N26626));
NAND2XL inst_cellmath__60_0_I527 (.Y(N3621), .A(N3593), .B(N3413));
NOR2XL inst_cellmath__60_0_I368 (.Y(N3402), .A(N3456), .B(N3446));
NOR2XL inst_cellmath__60_0_I348 (.Y(N3633), .A(N3603), .B(N3702));
ADDHX1 inst_cellmath__60_0_I16217 (.CO(N26603), .S(N26593), .A(N3402), .B(N3633));
ADDFX1 inst_cellmath__60_0_I16221 (.CO(N26590), .S(N26634), .A(N26603), .B(N26583), .CI(N26608));
AND2XL inst_cellmath__60_0_I16328 (.Y(N26636), .A(N26590), .B(N26596));
INVX1 inst_cellmath__60_0_I16240 (.Y(N26606), .A(N26634));
INVXL inst_cellmath__60_0_I377 (.Y(N3441), .A(N3412));
NOR2XL inst_cellmath__60_0_I347 (.Y(N3460), .A(N3603), .B(N3611));
ADDHX1 inst_cellmath__60_0_I16215 (.CO(N26610), .S(N3541), .A(N3441), .B(N3460));
NOR2XL inst_cellmath__60_0_I16214 (.Y(N26585), .A(N3503), .B(N3611));
ADDFX1 inst_cellmath__60_0_I16218 (.CO(N26629), .S(N26615), .A(N26610), .B(N26585), .CI(N26593));
INVXL inst_cellmath__60_0_I16239 (.Y(N26627), .A(N26629));
NAND2X1 inst_cellmath__60_0_I16237 (.Y(N26587), .A(N26629), .B(N26634));
INVX1 inst_cellmath__60_0_I16227 (.Y(N26616), .A(N26615));
NOR2XL inst_cellmath__60_0_I357 (.Y(N3623), .A(N3503), .B(N3446));
NOR2XL inst_cellmath__60_0_I367 (.Y(N3615), .A(N3456), .B(N3412));
NOR2XL inst_cellmath__60_0_I356 (.Y(N3452), .A(N3412), .B(N3503));
NOR2BX1 inst_cellmath__60_0_I346 (.Y(N3685), .AN(a_man[7]), .B(N3603));
ADDHXL inst_cellmath__60_0_I431 (.CO(N3451), .S(N3754), .A(N3452), .B(N3685));
ADDFXL inst_cellmath__60_0_I16216 (.CO(N26637), .S(N3712), .A(N3623), .B(N3615), .CI(N3451));
INVXL inst_cellmath__60_0_I16225 (.Y(N26624), .A(N26637));
NAND2X1 inst_cellmath__60_0_I16235 (.Y(N26638), .A(N26616), .B(N26624));
OR2XL inst_cellmath__60_0_I16329 (.Y(N26619), .A(N26624), .B(N26616));
AND2XL inst_cellmath__60_0_I492 (.Y(N3570), .A(N3541), .B(N3712));
INVXL inst_cellmath__60_0_I366 (.Y(N3668), .A(N3456));
NOR2BX1 inst_cellmath__60_0_I345 (.Y(N3511), .AN(a_man[6]), .B(N3603));
ADDHX1 inst_cellmath__60_0_I430 (.CO(N3673), .S(N3588), .A(N3668), .B(N3511));
NOR2XL inst_cellmath__60_0_I355 (.Y(N3674), .A(N3503), .B(N3456));
AND2XL inst_cellmath__60_0_I488 (.Y(N3617), .A(N3674), .B(N3588));
NOR3XL inst_cellmath__60_0_I5943 (.Y(N3555), .A(N3603), .B(N3503), .C(N3456));
OAI22XL inst_cellmath__60_0_I5861 (.Y(N3624), .A0(N3617), .A1(N3555), .B0(N3674), .B1(N3588));
NAND2XL inst_cellmath__60_0_I490 (.Y(N3404), .A(N3673), .B(N3754));
AOI2BB2X1 inst_cellmath__60_0_I5862 (.Y(N3526), .A0N(N3673), .A1N(N3754), .B0(N3624), .B1(N3404));
OAI22X1 inst_cellmath__60_0_I16234 (.Y(N26611), .A0(N3570), .A1(N3526), .B0(N3541), .B1(N3712));
OAI2BB1X1 inst_cellmath__60_0_I16282 (.Y(N26579), .A0N(N26619), .A1N(N26611), .B0(N26638));
AOI22X2 inst_cellmath__60_0_I16241 (.Y(N26581), .A0(N26627), .A1(N26606), .B0(N26587), .B1(N26579));
OR2XL inst_cellmath__60_0_I16285 (.Y(N26594), .A(N26590), .B(N26596));
OAI21X2 inst_cellmath__60_0_I16243 (.Y(N3753), .A0(N26636), .A1(N26581), .B0(N26594));
NOR2XL inst_cellmath__60_0_I526 (.Y(N3540), .A(N3593), .B(N3413));
AOI21X1 inst_cellmath__60_0_I554 (.Y(N3530), .A0(N3621), .A1(N3753), .B0(N3540));
NOR2X1 inst_cellmath__60_0_I528 (.Y(N3710), .A(N3489), .B(N3703));
NOR2XL inst_cellmath__60_0_I530 (.Y(N3483), .A(N3400), .B(N3771));
AOI21X2 inst_cellmath__60_0_I555 (.Y(N3475), .A0(N3574), .A1(N3710), .B0(N3483));
OAI21X1 inst_noninc_a_cellmath__55_2WWMM_I16169 (.Y(N3714), .A0(N3565), .A1(N3530), .B0(N3475));
NOR2X2 inst_noninc_a_cellmath__55_2WWMM_I16167 (.Y(N3657), .A(N3464), .B(N3619));
NOR2X1 inst_cellmath__60_0_I534 (.Y(N3438), .A(N3709), .B(N3694));
AOI21X4 inst_cellmath__60_0_I557 (.Y(N3430), .A0(N3657), .A1(N3521), .B0(N3438));
NOR2X2 inst_cellmath__60_0_I536 (.Y(N3605), .A(N3775), .B(N3590));
NOR2X1 inst_cellmath__60_0_I538 (.Y(N3392), .A(N3678), .B(N3486));
AOI21X4 inst_cellmath__60_0_I559 (.Y(N3768), .A0(N3605), .A1(N3471), .B0(N3392));
OAI21X2 inst_cellmath__60_0_I576 (.Y(N3662), .A0(N3463), .A1(N3430), .B0(N3768));
AOI21X1 inst_cellmath__60_0_I585 (.Y(N3509), .A0(N3714), .A1(N3742), .B0(N3662));
XNOR2XL inst_cellmath__60_0_I612 (.Y(inst_cellmath__60[17]), .A(N3491), .B(N3509));
INVX2 inst_cellmath__62_0_I1657 (.Y(N6446), .A(inst_cellmath__60[17]));
NOR2X1 inst_cellmath__62_0_I1787 (.Y(N6457), .A(N6347), .B(N6446));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1162 (.Y(N4385), .A(N4533), .B(N4413));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1163 (.Y(N4864), .A(N4385), .B(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I796 (.Y(N4692), .A(a_man[19]), .B(N4644));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1340 (.Y(N4543), .A(N4896), .B(N4692));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1554 (.Y(N4209), .A0(N4634), .A1(N4864), .B0(N4543), .B1(a_man[21]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1122 (.Y(N4867), .A(N4533), .B(N4349));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1123 (.Y(N4964), .A(N4867), .B(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1176 (.Y(N4563), .A(N4634), .B(N4964));
AO22XL inst_cellmath__62_0_I16290 (.Y(N6276), .A0(N4563), .A1(a_man[22]), .B0(N4911), .B1(N4209));
NOR2XL inst_cellmath__60_0_I418 (.Y(N3596), .A(N3432), .B(N3462));
INVXL inst_cellmath__60_0_I422 (.Y(N3569), .A(N3462));
NOR2XL inst_cellmath__60_0_I409 (.Y(N3537), .A(N3702), .B(N3538));
ADDFX1 inst_cellmath__60_0_I477 (.CO(N3474), .S(N3397), .A(N3596), .B(N3569), .CI(N3537));
OR2XL inst_cellmath__60_0_I403 (.Y(N3467), .A(N3611), .B(N3571));
NOR2XL inst_cellmath__60_0_I414 (.Y(N3453), .A(N3399), .B(N3496));
ADDFXL inst_cellmath__60_0_I478 (.CO(N3649), .S(N3564), .A(N3453), .B(N3467), .CI(N3743));
ADDFX1 inst_cellmath__60_0_I479 (.CO(N3429), .S(N3731), .A(N3529), .B(N3397), .CI(N3564));
NOR2XL inst_cellmath__60_0_I542 (.Y(N3726), .A(N3700), .B(N3731));
NAND2X1 inst_cellmath__60_0_I543 (.Y(N3426), .A(N3700), .B(N3731));
NAND2BXL inst_cellmath__60_0_I601 (.Y(N3747), .AN(N3726), .B(N3426));
XNOR2X1 inst_cellmath__60_0_I625 (.Y(N3696), .A(N3747), .B(N3642));
XNOR2X1 inst_cellmath__60_0_I626 (.Y(N3394), .A(N3747), .B(N3559));
MX2X1 inst_cellmath__62_0_I5908 (.Y(N6184), .A(N3696), .B(N3394), .S0(N3509));
NOR2X1 inst_cellmath__62_0_I1775 (.Y(N6392), .A(N6276), .B(N6184));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I745 (.Y(N5141), .A(a_man[17]), .B(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1457 (.Y(N4738), .A0(N4533), .A1(N5141), .B0(N5163), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I781 (.Y(N4633), .A(N4533), .B(N5141));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1504 (.Y(N4923), .A0(N4896), .A1(N4738), .B0(N4633), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1236 (.Y(N4261), .A(N4533), .B(N4849));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1339 (.Y(N4329), .A0(N4896), .A1(N4692), .B0(N4261), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1553 (.Y(N5006), .A0(N4634), .A1(N4923), .B0(N4329), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1077 (.Y(N4468), .A(N4619), .B(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1121 (.Y(N5093), .A(N4896), .B(N4468));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1175 (.Y(N4922), .A(a_man[21]), .B(N5093));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1606 (.Y(N456), .A0(N4911), .A1(N5006), .B0(N4922), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1756 (.Y(N6198), .A(N456));
NAND2X1 inst_cellmath__60_0_I562 (.Y(N3419), .A(N3426), .B(N3642));
NOR2X2 inst_cellmath__60_0_I579 (.Y(N3528), .A(N3419), .B(N3463));
NOR2X2 inst_cellmath__60_0_I575 (.Y(N3579), .A(N3565), .B(N3512));
NAND2X2 inst_cellmath__60_0_I587 (.Y(N3766), .A(N3528), .B(N3579));
INVXL inst_cellmath__60_0_I572 (.Y(N3589), .A(N3530));
INVXL inst_cellmath__60_0_I582 (.Y(N3675), .A(N3589));
OAI21X4 inst_cellmath__60_0_I574 (.Y(N3485), .A0(N3512), .A1(N3475), .B0(N3430));
AOI21X1 inst_cellmath__60_0_I561 (.Y(N3720), .A0(N3559), .A1(N3426), .B0(N3726));
OAI21X2 inst_cellmath__60_0_I578 (.Y(N3442), .A0(N3419), .A1(N3768), .B0(N3720));
AOI21X4 inst_cellmath__60_0_I586 (.Y(N3684), .A0(N3528), .A1(N3485), .B0(N3442));
OAI21X4 inst_noninc_a_cellmath__55_2WWMM_I16064 (.Y(N3534), .A0(N3766), .A1(N3675), .B0(N3684));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I16066 (.Y(N26104), .A(N3534));
NOR2XL inst_cellmath__60_0_I415 (.Y(N3625), .A(N3399), .B(N3538));
NOR2XL inst_cellmath__60_0_I419 (.Y(N3765), .A(N3432), .B(N3496));
OR2XL inst_cellmath__60_0_I410 (.Y(N3554), .A(N3702), .B(N3571));
ADDFX1 inst_cellmath__60_0_I480 (.CO(N3597), .S(N3510), .A(N3625), .B(N3765), .CI(N3554));
ADDFX1 inst_cellmath__60_0_I481 (.CO(N3767), .S(N3686), .A(N3510), .B(N3474), .CI(N3649));
NOR2XL inst_cellmath__60_0_I544 (.Y(N3504), .A(N3429), .B(N3686));
NAND2XL inst_cellmath__60_0_I545 (.Y(N3592), .A(N3429), .B(N3686));
NAND2BXL inst_noninc_a_cellmath__55_2WWMM_I16065 (.Y(N26096), .AN(N3504), .B(N3592));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I16067 (.Y(N26097), .A(N26096));
MXI2X1 inst_noninc_a_cellmath__55_2WWMM_I16071 (.Y(N26111), .A(N3534), .B(N26104), .S0(N26097));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I16076 (.Y(N6258), .A(N26111));
NOR2X2 inst_cellmath__62_0_I1763 (.Y(N6324), .A(N6198), .B(N6258));
ADDFHXL inst_cellmath__62_0_I1855 (.CO(N6493), .S(N6417), .A(N6457), .B(N6392), .CI(N6324));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1058 (.Y(N4584), .A0(N13806), .A1(N4166), .B0(N4736), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5884 (.Y(N5043), .A0(N4533), .A1(N4584), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5887 (.Y(N4648), .A0(N4896), .A1(N5043), .B0(N4852), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I879 (.Y(N4287), .A0(N4533), .A1(N5141), .B0(N5088), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I926 (.Y(N4683), .A0(N4896), .A1(N4287), .B0(N4633), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I16074 (.Y(N26095), .A0(N4634), .A1(N4648), .B0(N4683), .B1(a_man[21]));
NOR2X2 inst_noninc_a_cellmath__55_2WWMM_I677 (.Y(N4995), .A(N13760), .B(N13745));
CLKBUFX6 inst_noninc_a_cellmath__55_2WWMM_I5872 (.Y(N4297), .A(N4995));
NOR2X2 inst_noninc_a_cellmath__55_2WWMM_I6013 (.Y(N4438), .A(a_man[17]), .B(N13744));
AO22XL inst_noninc_a_cellmath__55_2WWMM_I821 (.Y(N5007), .A0(N13791), .A1(N4297), .B0(N4826), .B1(N4438));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I823 (.Y(N4162), .A(N5007));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1454 (.Y(N5094), .A0(N4533), .A1(N4162), .B0(N13745), .B1(a_man[19]));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5832 (.Y(N13797), .A(N13789));
NAND2X4 inst_noninc_a_cellmath__55_2WWMM_I734 (.Y(N4280), .A(N13744), .B(a_man[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I769 (.Y(N4377), .A0(N13797), .A1(N13744), .B0(N4280), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1398 (.Y(N5134), .A0(N4533), .A1(N4377), .B0(N4162), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1501 (.Y(N4255), .A0(N4896), .A1(N5094), .B0(N5134), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1053 (.Y(N4151), .A0(N13806), .A1(N13760), .B0(N4166), .B1(N13786));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I758 (.Y(N5061), .A0(N4826), .A1(N4479), .B0(N13791), .B1(a_man[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1233 (.Y(N4610), .A0(N4533), .A1(N4151), .B0(N5061), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1336 (.Y(N4677), .A0(N4896), .A1(N13766), .B0(N4610), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I16072 (.Y(N26089), .A0(N4634), .A1(N4255), .B0(N4677), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I16075 (.Y(N26100), .A0(a_man[22]), .A1(N26095), .B0(N26089), .B1(N4911));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I16077 (.Y(N6317), .A(N26100));
NOR2XL inst_cellmath__60_0_I427 (.Y(N3661), .A(N3496), .B(N3538));
INVXL inst_cellmath__60_0_I429 (.Y(N3683), .A(N3538));
OR2XL inst_cellmath__60_0_I425 (.Y(N3421), .A(N3462), .B(N3571));
ADDFX1 inst_cellmath__60_0_I485 (.CO(N3669), .S(N3584), .A(N3661), .B(N3683), .CI(N3421));
OR2XL inst_cellmath__60_0_I421 (.Y(N3724), .A(N3432), .B(N3571));
NOR2XL inst_cellmath__60_0_I424 (.Y(N3692), .A(N3462), .B(N3538));
NOR2XL inst_cellmath__60_0_I423 (.Y(N3518), .A(N3462), .B(N3496));
INVXL inst_cellmath__60_0_I426 (.Y(N3713), .A(N3496));
NOR2XL inst_cellmath__60_0_I420 (.Y(N3548), .A(N3432), .B(N3538));
ADDFX1 inst_cellmath__60_0_I482 (.CO(N3550), .S(N3461), .A(N3518), .B(N3713), .CI(N3548));
ADDFX1 inst_cellmath__60_0_I484 (.CO(N3494), .S(N3417), .A(N3724), .B(N3692), .CI(N3550));
NAND2XL inst_cellmath__60_0_I551 (.Y(N3717), .A(N3584), .B(N3494));
OR2XL inst_cellmath__60_0_I416 (.Y(N3637), .A(N3399), .B(N3571));
ADDFX1 inst_cellmath__60_0_I483 (.CO(N3719), .S(N3632), .A(N3597), .B(N3637), .CI(N3461));
NAND2XL inst_cellmath__60_0_I549 (.Y(N3545), .A(N3417), .B(N3719));
NAND2XL inst_cellmath__60_0_I568 (.Y(N3708), .A(N3717), .B(N3545));
NAND2XL inst_cellmath__60_0_I547 (.Y(N3760), .A(N3767), .B(N3632));
NAND2XL inst_cellmath__60_0_I564 (.Y(N3751), .A(N3760), .B(N3592));
OR2XL inst_cellmath__60_0_I571 (.Y(N3500), .A(N3751), .B(N3708));
NOR2XL inst_cellmath__60_0_I581 (.Y(N3699), .A(N3419), .B(N3500));
NAND2XL inst_cellmath__60_0_I589 (.Y(N3549), .A(N3699), .B(N3742));
INVXL inst_noninc_a_cellmath__55_2WWMM_I16170 (.Y(N3756), .A(N3714));
NOR2XL inst_cellmath__60_0_I546 (.Y(N3679), .A(N3767), .B(N3632));
AOI21XL inst_cellmath__60_0_I563 (.Y(N3670), .A0(N3760), .A1(N3504), .B0(N3679));
NOR2XL inst_cellmath__60_0_I548 (.Y(N3455), .A(N3417), .B(N3719));
NOR2XL inst_cellmath__60_0_I550 (.Y(N3627), .A(N3584), .B(N3494));
AOI21XL inst_cellmath__60_0_I567 (.Y(N3618), .A0(N3717), .A1(N3455), .B0(N3627));
OA21X1 inst_cellmath__60_0_I570 (.Y(N3424), .A0(N3708), .A1(N3670), .B0(N3618));
OAI21X1 inst_cellmath__60_0_I580 (.Y(N3608), .A0(N3500), .A1(N3720), .B0(N3424));
AOI21XL inst_cellmath__60_0_I588 (.Y(N3459), .A0(N3699), .A1(N3662), .B0(N3608));
OAI21X1 inst_cellmath__60_0_I591 (.Y(N3705), .A0(N3549), .A1(N3756), .B0(N3459));
OR2XL inst_cellmath__60_0_I428 (.Y(N3499), .A(N3496), .B(N3571));
NOR2XL inst_cellmath__60_0_I552 (.Y(N3411), .A(N3499), .B(N3669));
NAND2XL inst_cellmath__60_0_I553 (.Y(N3488), .A(N3499), .B(N3669));
NAND2BXL inst_cellmath__60_0_I606 (.Y(N3466), .AN(N3411), .B(N3488));
XNOR2X1 inst_cellmath__62_0_I5913 (.Y(N6213), .A(N3705), .B(N3466));
NOR2XL inst_cellmath__62_0_I1728 (.Y(N6274), .A(N6317), .B(N6213));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I645 (.Y(N4206), .A(N13745));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5783 (.Y(N13748), .A(N4206));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5789 (.Y(N13754), .A(N13748));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I845 (.Y(N4939), .A0(N13803), .A1(N4736), .B0(N13754), .B1(N13782));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I735 (.Y(N4713), .A0(N13760), .A1(N13744), .B0(N13745), .B1(a_man[17]));
CLKINVX4 inst_noninc_a_cellmath__55_2WWMM_I736 (.Y(N5081), .A(N4713));
INVX12 inst_noninc_a_cellmath__55_2WWMM_I737 (.Y(N4953), .A(N5081));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I992 (.Y(N4820), .A(N13795), .B(N4953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1452 (.Y(N4649), .A0(N4533), .A1(N4939), .B0(N4820), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I839 (.Y(N4435), .A0(N13745), .A1(N4826), .B0(N13803), .B1(N4953));
NAND2X4 inst_noninc_a_cellmath__55_2WWMM_I665 (.Y(N4300), .A(N13745), .B(N13760));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1002 (.Y(N4207), .A0(N13786), .A1(N4300), .B0(N13795), .B1(N13745));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1396 (.Y(N4682), .A0(N4533), .A1(N4435), .B0(N4207), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1499 (.Y(N4829), .A0(N4896), .A1(N4649), .B0(N4682), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1293 (.Y(N4632), .A0(N4533), .A1(N4349), .B0(N5088), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I708 (.Y(N4929), .A0(N4314), .A1(N4869), .B0(a_man[17]), .B1(N4826));
AOI22X4 inst_noninc_a_cellmath__55_2WWMM_I746 (.Y(N4457), .A0(N13795), .A1(N4953), .B0(N4280), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1231 (.Y(N4165), .A0(N4533), .A1(N4929), .B0(N4457), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1334 (.Y(N4234), .A0(N4896), .A1(N4632), .B0(N4165), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1548 (.Y(N4919), .A0(N4634), .A1(N4829), .B0(N4234), .B1(a_man[21]));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5787 (.Y(N13752), .A(N13748));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1057 (.Y(N4268), .A0(N13806), .A1(N4953), .B0(N13752), .B1(N13786));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I5883 (.Y(N4875), .A0(N4206), .A1(N4314), .B0(N4300), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1073 (.Y(N4597), .A0(N4533), .A1(N4268), .B0(N4875), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I850 (.Y(N4805), .A0(N13803), .A1(N13745), .B0(N4297), .B1(N13782));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5807 (.Y(N13772), .A(N13767));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I968 (.Y(N4783), .A0(N4280), .A1(N13803), .B0(N4300), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1005 (.Y(N4323), .A0(N4533), .A1(N4805), .B0(N4783), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1117 (.Y(N4203), .A0(N4896), .A1(N4597), .B0(N4323), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I830 (.Y(N4879), .A0(N13797), .A1(N4953), .B0(N13760), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I877 (.Y(N4857), .A0(N4533), .A1(N4879), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I710 (.Y(N5078), .A0(N4314), .A1(N4166), .B0(N4869), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I779 (.Y(N4186), .A0(a_man[17]), .A1(N4533), .B0(N5078), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I924 (.Y(N4240), .A0(N4896), .A1(N4857), .B0(N4186), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1169 (.Y(N4605), .A0(N4634), .A1(N4203), .B0(N4240), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1601 (.Y(N451), .A0(N4911), .A1(N4919), .B0(N4605), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1691 (.Y(N6509), .A(N451));
NOR2BX1 inst_cellmath__60_0_I607 (.Y(N3723), .AN(N3538), .B(N3571));
XNOR2X1 inst_cellmath__60_0_I641 (.Y(N3629), .A(N3723), .B(N3411));
XNOR2X1 inst_cellmath__60_0_I640 (.Y(N3546), .A(N3723), .B(N3488));
MX2X1 inst_cellmath__62_0_I5914 (.Y(N6286), .A(N3629), .B(N3546), .S0(N3705));
NOR2X1 inst_cellmath__62_0_I1703 (.Y(N6330), .A(N6509), .B(N6286));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I16172 (.Y(N26412), .A(N4634), .B(N5093));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I754 (.Y(N4768), .A0(N4869), .A1(N13791), .B0(N4826), .B1(N4479));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1456 (.Y(N4515), .A0(N4344), .A1(N4533), .B0(a_man[19]), .B1(N4768));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I855 (.Y(N4674), .A0(N13806), .A1(N4869), .B0(N13760), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1400 (.Y(N4547), .A0(N4533), .A1(N4674), .B0(N4349), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1503 (.Y(N4694), .A0(N4896), .A1(N4515), .B0(N4547), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1295 (.Y(N4720), .A0(N4533), .A1(N4644), .B0(N4968), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1235 (.Y(N5055), .A0(N4533), .A1(N4341), .B0(N4413), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1338 (.Y(N5128), .A0(N4896), .A1(N4720), .B0(N5055), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I16173 (.Y(N26419), .A0(N4634), .A1(N4694), .B0(N5128), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I16175 (.Y(N26399), .A0(N26412), .A1(a_man[22]), .B0(N4911), .B1(N26419));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I16176 (.Y(N6467), .A(N26399));
NAND2BXL inst_cellmath__60_0_I603 (.Y(N3478), .AN(N3679), .B(N3760));
XNOR2X1 inst_cellmath__60_0_I629 (.Y(N3644), .A(N3478), .B(N3504));
XNOR2X1 inst_cellmath__60_0_I628 (.Y(N3560), .A(N3478), .B(N3592));
MX2X1 inst_cellmath__62_0_I5910 (.Y(N6331), .A(N3644), .B(N3560), .S0(N3534));
NOR2XL inst_cellmath__62_0_I1751 (.Y(N6260), .A(N6467), .B(N6331));
NAND2BXL inst_cellmath__60_0_I605 (.Y(N3600), .AN(N3627), .B(N3717));
INVXL inst_cellmath__60_0_I566 (.Y(N3480), .A(N3545));
INVXL inst_cellmath__60_0_I565 (.Y(N3403), .A(N3455));
OAI21XL inst_cellmath__60_0_I569 (.Y(N3737), .A0(N3480), .A1(N3670), .B0(N3403));
XNOR2X1 inst_cellmath__60_0_I635 (.Y(N3680), .A(N3600), .B(N3737));
NOR2XL inst_cellmath__60_0_I636 (.Y(N3704), .A(N3480), .B(N3751));
NOR2XL inst_cellmath__60_0_I637 (.Y(N3582), .A(N3704), .B(N3737));
XOR2XL inst_cellmath__60_0_I638 (.Y(N3762), .A(N3600), .B(N3582));
MX2X1 inst_cellmath__62_0_I5912 (.Y(N6477), .A(N3680), .B(N3762), .S0(N3534));
NOR2XL inst_cellmath__62_0_I1727 (.Y(N6465), .A(N6317), .B(N6477));
ADDFXL inst_cellmath__62_0_I1856 (.CO(N6299), .S(N6228), .A(N6330), .B(N6260), .CI(N6465));
ADDFX1 inst_cellmath__62_0_I1864 (.CO(N6468), .S(N6394), .A(N6493), .B(N6274), .CI(N6299));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I841 (.Y(N5108), .A0(N4826), .A1(N4953), .B0(N4300), .B1(N13803));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1453 (.Y(N4872), .A0(N4533), .A1(N5108), .B0(N4349), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1050 (.Y(N4392), .A0(N13806), .A1(N4479), .B0(N4953), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1397 (.Y(N4907), .A0(N4533), .A1(N4392), .B0(N4457), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1500 (.Y(N5050), .A0(N4896), .A1(N4872), .B0(N4907), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1222 (.Y(N4951), .A0(N4314), .A1(N4280), .B0(N4953), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1232 (.Y(N4386), .A0(N4533), .A1(N4951), .B0(N4783), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1335 (.Y(N4455), .A0(N4896), .A1(N13754), .B0(N4386), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1549 (.Y(N5142), .A0(N4634), .A1(N5050), .B0(N4455), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I862 (.Y(N4540), .A0(N13806), .A1(N4297), .B0(N13782), .B1(N4953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1047 (.Y(N5046), .A0(N13795), .A1(N4953), .B0(N4869), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1074 (.Y(N4819), .A0(N4533), .A1(N4540), .B0(N5046), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I981 (.Y(N4786), .A0(N13795), .A1(a_man[17]), .B0(N4736), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1006 (.Y(N4538), .A0(N4786), .A1(N4533), .B0(a_man[19]), .B1(N4276));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1118 (.Y(N4422), .A0(N4896), .A1(N4819), .B0(N4538), .B1(a_man[20]));
XNOR2X1 inst_noninc_a_cellmath__55_2WWMM_I6016 (.Y(N4469), .A(N4826), .B(a_man[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I878 (.Y(N5079), .A0(N4533), .A1(N4344), .B0(N4469), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I780 (.Y(N4408), .A0(N4533), .A1(N4469), .B0(N4349), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I925 (.Y(N4463), .A0(N4896), .A1(N5079), .B0(N4408), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1171 (.Y(N4828), .A0(N4634), .A1(N4422), .B0(N4463), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1602 (.Y(N452), .A0(N4911), .A1(N5142), .B0(N4828), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1704 (.Y(N6244), .A(N452));
NOR2X1 inst_cellmath__62_0_I1714 (.Y(N6251), .A(N6244), .B(N6477));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I859 (.Y(N5159), .A(N13806), .B(N4280));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1388 (.Y(N5087), .A0(N4314), .A1(N13754), .B0(N4438), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1451 (.Y(N4423), .A0(N4533), .A1(N5159), .B0(N5087), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I984 (.Y(N4774), .A0(N13745), .A1(N13795), .B0(a_man[17]), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1001 (.Y(N5062), .A0(N13795), .A1(N13760), .B0(N4280), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1395 (.Y(N4462), .A0(N4533), .A1(N4774), .B0(N5062), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1498 (.Y(N4606), .A0(N4896), .A1(N4423), .B0(N4462), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I999 (.Y(N4519), .A(N13806), .B(a_man[17]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1292 (.Y(N4407), .A0(N4533), .A1(N5046), .B0(N4519), .B1(a_man[19]));
INVX2 inst_noninc_a_cellmath__55_2WWMM_I5798 (.Y(N13763), .A(N13761));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I840 (.Y(N4948), .A0(N4280), .A1(N13803), .B0(N13763), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1230 (.Y(N4963), .A0(N4533), .A1(N4268), .B0(N4948), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1333 (.Y(N5031), .A0(N4896), .A1(N4407), .B0(N4963), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1547 (.Y(N4690), .A0(N4634), .A1(N4606), .B0(N5031), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1042 (.Y(N4372), .A(N4736), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1072 (.Y(N4370), .A0(N4533), .A1(N4341), .B0(N4372), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I861 (.Y(N5124), .A0(N13806), .A1(N13760), .B0(N4953), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1004 (.Y(N5120), .A0(N4533), .A1(N5124), .B0(N4457), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1116 (.Y(N5000), .A0(N4896), .A1(N4370), .B0(N5120), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I853 (.Y(N4307), .A0(N13803), .A1(N13754), .B0(N13745), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I876 (.Y(N4637), .A0(N4533), .A1(N4307), .B0(N13752), .B1(a_man[19]));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5797 (.Y(N13762), .A(N13761));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I709 (.Y(N4856), .A0(N4314), .A1(N4995), .B0(N13762), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I778 (.Y(N4983), .A0(N4533), .A1(N13752), .B0(N4856), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I923 (.Y(N5037), .A0(N4896), .A1(N4637), .B0(N4983), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1168 (.Y(N4379), .A0(N4634), .A1(N5000), .B0(N5037), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1600 (.Y(N450), .A0(N4911), .A1(N4690), .B0(N4379), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1678 (.Y(N6434), .A(N450));
NOR2X1 inst_cellmath__62_0_I1690 (.Y(N6452), .A(N6434), .B(N6286));
NAND2BXL inst_cellmath__60_0_I604 (.Y(N3734), .AN(N3455), .B(N3545));
INVXL inst_cellmath__60_0_I592 (.Y(N3647), .A(N3670));
XNOR2X1 inst_cellmath__60_0_I631 (.Y(N3427), .A(N3734), .B(N3647));
NOR2BX1 inst_cellmath__60_0_I632 (.Y(N3594), .AN(N3751), .B(N3647));
XOR2XL inst_cellmath__60_0_I633 (.Y(N3506), .A(N3734), .B(N3594));
MX2X1 inst_cellmath__62_0_I5911 (.Y(N6404), .A(N3427), .B(N3506), .S0(N3534));
NOR2XL inst_cellmath__62_0_I1726 (.Y(N6316), .A(N6317), .B(N6404));
ADDFX1 inst_cellmath__62_0_I1849 (.CO(N6285), .S(N6209), .A(N6452), .B(N6251), .CI(N6316));
NOR2X1 inst_cellmath__62_0_I1750 (.Y(N6449), .A(N6467), .B(N6258));
NOR2XL inst_cellmath__62_0_I1762 (.Y(N6178), .A(N6198), .B(N6184));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1455 (.Y(N4301), .A0(N4533), .A1(N4457), .B0(N4739), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I990 (.Y(N5101), .A0(N13795), .A1(N13763), .B0(N13760), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1399 (.Y(N4335), .A0(N4533), .A1(N5101), .B0(N4706), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1502 (.Y(N4476), .A0(N4896), .A1(N4301), .B0(N4335), .B1(a_man[20]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I1294 (.Y(N4503), .A(N4252));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1234 (.Y(N4834), .A0(N4533), .A1(N4271), .B0(N5163), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1337 (.Y(N4901), .A0(N4896), .A1(N4503), .B0(N4834), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1551 (.Y(N4559), .A0(N4634), .A1(N4476), .B0(N4901), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5885 (.Y(N4247), .A0(N4533), .A1(N4349), .B0(N4619), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I917 (.Y(N4718), .A(N4533), .B(N13803));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5888 (.Y(N4871), .A0(N4896), .A1(N4247), .B0(N4718), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I880 (.Y(N4505), .A(N4533), .B(N5141));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I927 (.Y(N4908), .A(a_man[20]), .B(N4505));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5892 (.Y(N4254), .A0(N4634), .A1(N4871), .B0(N4908), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1604 (.Y(N454), .A0(N4911), .A1(N4559), .B0(N4254), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1730 (.Y(N6391), .A(N454));
NOR2XL inst_cellmath__62_0_I1738 (.Y(N6381), .A(N6391), .B(N6331));
ADDFXL inst_cellmath__62_0_I1848 (.CO(N6474), .S(N6401), .A(N6449), .B(N6178), .CI(N6381));
ADDFHXL inst_cellmath__62_0_I1858 (.CO(N6259), .S(N6185), .A(N6285), .B(N6474), .CI(N6417));
NOR2XL inst_cellmath__62_0_I1702 (.Y(N6183), .A(N6509), .B(N6213));
NOR2X2 inst_cellmath__62_0_I1774 (.Y(N6245), .A(N6276), .B(N6446));
NAND2BXL inst_cellmath__60_0_I599 (.Y(N3631), .AN(N3392), .B(N3471));
XNOR2XL inst_cellmath__60_0_I622 (.Y(N3439), .A(N3695), .B(N3631));
XNOR2XL inst_cellmath__60_0_I623 (.Y(N3523), .A(N3605), .B(N3631));
AOI21X2 inst_cellmath__60_0_I584 (.Y(N3730), .A0(N3579), .A1(N3589), .B0(N3485));
MX2X1 inst_cellmath__62_0_I5906 (.Y(N6372), .A(N3439), .B(N3523), .S0(N3730));
NOR2X1 inst_cellmath__62_0_I1786 (.Y(N6310), .A(N6347), .B(N6372));
ADDHX1 inst_cellmath__62_0_I1847 (.CO(N6327), .S(N6255), .A(N6245), .B(N6310));
NOR2XL inst_cellmath__62_0_I1749 (.Y(N6301), .A(N6467), .B(N6184));
NOR2X1 inst_cellmath__62_0_I1773 (.Y(N6435), .A(N6276), .B(N6372));
NOR2X1 inst_cellmath__62_0_I1761 (.Y(N6367), .A(N6198), .B(N6446));
ADDFXL inst_cellmath__62_0_I1839 (.CO(N6499), .S(N6423), .A(N6367), .B(N6435), .CI(N6301));
ADDFXL inst_cellmath__62_0_I1850 (.CO(N6431), .S(N6357), .A(N6255), .B(N6183), .CI(N6499));
NOR2X1 inst_cellmath__62_0_I1739 (.Y(N6191), .A(N6391), .B(N6404));
NOR2XL inst_cellmath__62_0_I1715 (.Y(N6397), .A(N6244), .B(N6213));
ADDFXL inst_cellmath__62_0_I1857 (.CO(N6447), .S(N6374), .A(N6191), .B(N6327), .CI(N6397));
ADDFX1 inst_cellmath__62_0_I1859 (.CO(N6405), .S(N6333), .A(N6431), .B(N6228), .CI(N6374));
ADDFHXL inst_cellmath__62_0_I1866 (.CO(N6422), .S(N6350), .A(N6394), .B(N6259), .CI(N6405));
NOR2XL inst_cellmath__62_0_I1740 (.Y(N6342), .A(N6391), .B(N6477));
NOR2X1 inst_cellmath__62_0_I1716 (.Y(N6204), .A(N6244), .B(N6286));
NOR2XL inst_cellmath__62_0_I1752 (.Y(N6407), .A(N6467), .B(N6404));
ADDFXL inst_cellmath__62_0_I1863 (.CO(N6318), .S(N6247), .A(N6204), .B(N6342), .CI(N6407));
NOR2X1 inst_cellmath__62_0_I1776 (.Y(N6199), .A(N6276), .B(N6258));
NOR2XL inst_cellmath__62_0_I1788 (.Y(N6269), .A(N6347), .B(N6184));
NOR2XL inst_cellmath__62_0_I1764 (.Y(N6473), .A(N6198), .B(N6331));
ADDFXL inst_cellmath__62_0_I1862 (.CO(N6510), .S(N6436), .A(N6199), .B(N6269), .CI(N6473));
NOR2XL inst_cellmath__62_0_I1777 (.Y(N6348), .A(N6276), .B(N6331));
NOR2XL inst_cellmath__62_0_I1789 (.Y(N6415), .A(N6347), .B(N6258));
NOR2XL inst_cellmath__62_0_I1729 (.Y(N6420), .A(N6317), .B(N6286));
ADDFX1 inst_cellmath__62_0_I1868 (.CO(N6379), .S(N6306), .A(N6348), .B(N6415), .CI(N6420));
ADDFX1 inst_cellmath__62_0_I1870 (.CO(N6339), .S(N6265), .A(N6318), .B(N6510), .CI(N6306));
NOR2XL inst_cellmath__62_0_I1765 (.Y(N6283), .A(N6198), .B(N6404));
NOR2XL inst_cellmath__62_0_I1753 (.Y(N6216), .A(N6467), .B(N6477));
NOR2XL inst_cellmath__62_0_I1741 (.Y(N6489), .A(N6391), .B(N6213));
ADDFX1 inst_cellmath__62_0_I1869 (.CO(N6189), .S(N6453), .A(N6283), .B(N6216), .CI(N6489));
ADDFXL inst_cellmath__62_0_I1865 (.CO(N6277), .S(N6200), .A(N6447), .B(N6436), .CI(N6247));
ADDFXL inst_cellmath__62_0_I1871 (.CO(N6486), .S(N6409), .A(N6468), .B(N6453), .CI(N6277));
ADDFHXL inst_cellmath__62_0_I1872 (.CO(inst_cellmath__62__W0[20]), .S(inst_cellmath__62__W1[19]), .A(N6422), .B(N6265), .CI(N6409));
NOR2XL inst_cellmath__62_0_I1701 (.Y(N6373), .A(N6509), .B(N6477));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I973 (.Y(N4704), .A(N13791), .B(N4953));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I725 (.Y(N4531), .A0(N4314), .A1(N4166), .B0(N4300), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1450 (.Y(N4204), .A0(N4533), .A1(N4704), .B0(N4531), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1066 (.Y(N4270), .A0(N13807), .A1(N4297), .B0(N4479), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1394 (.Y(N4239), .A0(N4533), .A1(N4162), .B0(N4270), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1497 (.Y(N4380), .A0(N4896), .A1(N4204), .B0(N4239), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I860 (.Y(N4897), .A0(N13806), .A1(N13760), .B0(N13754), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1291 (.Y(N4185), .A0(N4533), .A1(N4856), .B0(N4897), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1055 (.Y(N5140), .A0(N13806), .A1(N4438), .B0(N13752), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1229 (.Y(N4735), .A0(N4533), .A1(N4341), .B0(N5140), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1332 (.Y(N4809), .A0(N4896), .A1(N4185), .B0(N4735), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1546 (.Y(N4472), .A0(N4634), .A1(N4380), .B0(N4809), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1056 (.Y(N4496), .A0(N13806), .A1(N4438), .B0(N4869), .B1(N13786));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I874 (.Y(N4290), .A(N13803), .B(N4736));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1071 (.Y(N4153), .A0(N4533), .A1(N4496), .B0(N4290), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I976 (.Y(N4471), .A0(N13791), .A1(N4300), .B0(N13745), .B1(N13782));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I967 (.Y(N4154), .A0(N13803), .A1(N4438), .B0(N4300), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1003 (.Y(N4892), .A0(N4533), .A1(N4471), .B0(N4154), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1115 (.Y(N4776), .A0(N4896), .A1(N4153), .B0(N4892), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I761 (.Y(N5004), .A(N13795), .B(a_man[17]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I875 (.Y(N4189), .A(N4533), .B(N5004));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I777 (.Y(N4758), .A0(N4533), .A1(N5163), .B0(N4929), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I921 (.Y(N4814), .A0(N4896), .A1(N4189), .B0(N4758), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1167 (.Y(N4161), .A0(N4634), .A1(N4776), .B0(N4814), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1599 (.Y(N449), .A0(N4911), .A1(N4472), .B0(N4161), .B1(a_man[22]));
INVX1 inst_cellmath__62_0_I1665 (.Y(N6359), .A(N449));
NOR2XL inst_cellmath__62_0_I1677 (.Y(N6239), .A(N6359), .B(N6286));
NOR2XL inst_cellmath__62_0_I1713 (.Y(N6440), .A(N6244), .B(N6404));
ADDFX1 inst_cellmath__62_0_I1841 (.CO(N6455), .S(N6380), .A(N6373), .B(N6239), .CI(N6440));
NOR2XL inst_cellmath__62_0_I1737 (.Y(N6234), .A(N6391), .B(N6258));
NAND2BXL inst_cellmath__60_0_I598 (.Y(N3763), .AN(N3605), .B(N3695));
CLKXOR2X1 inst_cellmath__62_0_I5905 (.Y(N6298), .A(N3730), .B(N3763));
NOR2XL inst_cellmath__62_0_I1785 (.Y(N6501), .A(N6347), .B(N6298));
NOR2XL inst_cellmath__62_0_I1725 (.Y(N6508), .A(N6317), .B(N6331));
ADDFXL inst_cellmath__62_0_I1840 (.CO(N6308), .S(N6233), .A(N6501), .B(N6508), .CI(N6234));
ADDFXL inst_cellmath__62_0_I1851 (.CO(N6238), .S(N6505), .A(N6455), .B(N6308), .CI(N6401));
NAND2BXL inst_cellmath__60_0_I597 (.Y(N3508), .AN(N3438), .B(N3521));
XNOR2X1 inst_cellmath__60_0_I619 (.Y(N3575), .A(N3739), .B(N3508));
XNOR2X1 inst_cellmath__60_0_I620 (.Y(N3659), .A(N3657), .B(N3508));
MX2X1 inst_cellmath__62_0_I5904 (.Y(N6227), .A(N3575), .B(N3659), .S0(N3756));
NOR2X1 inst_cellmath__62_0_I1784 (.Y(N6353), .A(N6347), .B(N6227));
NOR2X1 inst_cellmath__62_0_I1736 (.Y(N6424), .A(N6391), .B(N6184));
NOR2XL inst_cellmath__62_0_I1760 (.Y(N6220), .A(N6198), .B(N6372));
ADDFXL inst_cellmath__62_0_I1831 (.CO(N6336), .S(N6262), .A(N6353), .B(N6424), .CI(N6220));
NOR2XL inst_cellmath__62_0_I1689 (.Y(N6307), .A(N6434), .B(N6213));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I16294 (.Y(N26090), .A(N3534), .B(N26096));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I16068 (.Y(N26108), .A(N26097), .B(N26104));
NOR3X1 inst_noninc_a_cellmath__55_2WWMM_I16078 (.Y(N6358), .A(N6317), .B(N26090), .C(N26108));
NOR2XL inst_cellmath__62_0_I1748 (.Y(N6494), .A(N6467), .B(N6446));
NOR2XL inst_cellmath__62_0_I1772 (.Y(N6287), .A(N6276), .B(N6298));
ADDFX1 inst_cellmath__62_0_I1832 (.CO(N6482), .S(N6408), .A(N6494), .B(N6358), .CI(N6287));
ADDFXL inst_cellmath__62_0_I1842 (.CO(N6267), .S(N6190), .A(N6307), .B(N6336), .CI(N6482));
ADDFXL inst_cellmath__64_0_I16106 (.CO(N6386), .S(N26219), .A(N6267), .B(N6209), .CI(N6357));
ADDFHXL inst_cellmath__62_0_I1860 (.CO(N6214), .S(N6480), .A(N6238), .B(N6185), .CI(N6386));
ADDFXL inst_cellmath__62_0_I1867 (.CO(inst_cellmath__62__W0[19]), .S(inst_cellmath__62__W1[18]), .A(N6214), .B(N6200), .CI(N6350));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1091 (.Y(N4705), .A0(N4533), .A1(N4849), .B0(N4644), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1020 (.Y(N5001), .A0(N4533), .A1(N4968), .B0(N4341), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1137 (.Y(N4888), .A0(N4896), .A1(N4705), .B0(a_man[20]), .B1(N5001));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I894 (.Y(N4726), .A(N4533), .B(N4413));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I941 (.Y(N4925), .A0(N4896), .A1(N4726), .B0(N4692), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1190 (.Y(N5068), .A0(N4888), .A1(N4634), .B0(N4925), .B1(a_man[21]));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I975 (.Y(N5045), .A0(N13791), .A1(N4953), .B0(a_man[17]), .B1(N13772));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1471 (.Y(N5116), .A0(N4533), .A1(a_man[17]), .B0(a_man[19]), .B1(N5045));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1391 (.Y(N5096), .A0(N4314), .A1(N4479), .B0(N4166), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1414 (.Y(N4695), .A0(N4533), .A1(N5096), .B0(a_man[19]), .B1(N4469));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1518 (.Y(N4844), .A0(N4896), .A1(N5116), .B0(a_man[20]), .B1(N4695));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I893 (.Y(N4873), .A0(N4533), .A1(N4413), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1354 (.Y(N4473), .A0(N4896), .A1(N4408), .B0(N4873), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1570 (.Y(N4936), .A0(N4634), .A1(N4844), .B0(N4473), .B1(a_man[21]));
AOI22X1 inst_cellmath__63_0_I5921 (.Y(N7645), .A0(N5068), .A1(a_man[22]), .B0(N4911), .B1(N4936));
INVX2 inst_cellmath__63_0_I1914 (.Y(N6952), .A(N7645));
NOR2XL inst_cellmath__63_0_I1973 (.Y(N6852), .A(N3142), .B(N6952));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1447 (.Y(N4916), .A(N13782), .B(N13766));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I765 (.Y(N4740), .A0(N13797), .A1(N4297), .B0(N4280), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1465 (.Y(N4797), .A0(N4916), .A1(N4533), .B0(a_man[19]), .B1(N4740));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1069 (.Y(N4357), .A(N13786), .B(N13752));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I764 (.Y(N4517), .A0(a_man[17]), .A1(N13797), .B0(N4297), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1408 (.Y(N4381), .A0(N4357), .A1(N4533), .B0(N4517), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1512 (.Y(N4525), .A0(N4896), .A1(N4797), .B0(N4381), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I972 (.Y(N4489), .A0(N13803), .A1(N4736), .B0(N4280), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1273 (.Y(N4912), .A0(N4314), .A1(N13760), .B0(N4300), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1303 (.Y(N4201), .A0(N4533), .A1(N4489), .B0(N4912), .B1(a_man[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1224 (.Y(N5098), .A(N4314), .B(N13754));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1244 (.Y(N4887), .A0(N4533), .A1(N5098), .B0(N4341), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1348 (.Y(N4157), .A0(N4896), .A1(N4201), .B0(N4887), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1564 (.Y(N4617), .A0(N4634), .A1(N4525), .B0(N4157), .B1(a_man[21]));
AO22XL inst_noninc_a_cellmath__55_2WWMM_I770 (.Y(N4825), .A0(N4613), .A1(N4314), .B0(N4300), .B1(N4826));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I772 (.Y(N5022), .A(N4825));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1085 (.Y(N4742), .A0(N4533), .A1(N5022), .B0(N4372), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1014 (.Y(N4688), .A0(N13745), .A1(N4533), .B0(a_man[19]), .B1(N4276));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1131 (.Y(N4569), .A0(N4896), .A1(N4742), .B0(a_man[20]), .B1(N4688));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I829 (.Y(N4431), .A0(N13797), .A1(N13745), .B0(N13754), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I888 (.Y(N4780), .A0(N4533), .A1(N5124), .B0(a_man[19]), .B1(N4431));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I751 (.Y(N4903), .A0(N13745), .A1(N13795), .B0(N13762), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I789 (.Y(N4910), .A0(N4533), .A1(N4903), .B0(N4271), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I935 (.Y(N4608), .A0(N4896), .A1(N4780), .B0(a_man[20]), .B1(N4910));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1184 (.Y(N4749), .A0(N4634), .A1(N4569), .B0(a_man[21]), .B1(N4608));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1616 (.Y(inst_cellmath__51[7]), .A0(N4617), .A1(N4911), .B0(a_man[22]), .B1(N4749));
INVX2 inst_cellmath__63_0_I1902 (.Y(N7016), .A(inst_cellmath__51[7]));
NOR2XL inst_cellmath__63_0_I2081 (.Y(N7029), .A(N3611), .B(N7016));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1470 (.Y(N4889), .A0(N4875), .A1(N4533), .B0(a_man[19]), .B1(N4431));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I5727 (.Y(N13558), .A0(N13791), .A1(N4438), .B0(N13788), .B1(N13762));
BUFX3 inst_noninc_a_cellmath__55_2WWMM_I5881 (.Y(N4177), .A(N13558));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1062 (.Y(N4745), .A0(N4300), .A1(N13807), .B0(a_man[17]), .B1(N13786));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1413 (.Y(N4477), .A0(N4533), .A1(N4177), .B0(a_man[19]), .B1(N4745));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1517 (.Y(N4622), .A0(N4896), .A1(N4889), .B0(a_man[20]), .B1(N4477));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I768 (.Y(N4615), .A0(N13797), .A1(N4736), .B0(N4479), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1308 (.Y(N4298), .A0(N4533), .A1(N13760), .B0(N4615), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1353 (.Y(N4251), .A0(N4298), .A1(N4896), .B0(a_man[20]), .B1(N4651));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1569 (.Y(N4707), .A0(N4634), .A1(N4622), .B0(a_man[21]), .B1(N4251));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1090 (.Y(N4490), .A0(N4533), .A1(N5061), .B0(a_man[19]), .B1(N4768));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I977 (.Y(N4918), .A0(N13791), .A1(a_man[17]), .B0(N4166), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1019 (.Y(N4778), .A0(N4533), .A1(N4674), .B0(N4918), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1136 (.Y(N4667), .A0(N4896), .A1(N4490), .B0(N4778), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I795 (.Y(N4997), .A(a_man[19]), .B(N4968));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I940 (.Y(N4696), .A0(N4873), .A1(N4896), .B0(N4997), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1189 (.Y(N4843), .A0(N4634), .A1(N4667), .B0(a_man[21]), .B1(N4696));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1621 (.Y(inst_cellmath__51[12]), .A0(N4911), .A1(N4707), .B0(N4843), .B1(a_man[22]));
CLKBUFX2 inst_cellmath__63_0_I1911 (.Y(N7067), .A(inst_cellmath__51[12]));
INVX3 inst_cellmath__63_0_I1912 (.Y(N7257), .A(N7067));
NOR2XL inst_cellmath__63_0_I1991 (.Y(N6880), .A(N3603), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2320 (.CO(N7614), .S(N7421), .A(N7029), .B(N6852), .CI(N6880));
INVX1 inst_cellmath__63_0_I1940 (.Y(N7350), .A(a_man[1]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1092 (.Y(N4934), .A(a_man[19]), .B(N4341));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1138 (.Y(N5115), .A0(N4896), .A1(N4934), .B0(N4279), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I813 (.Y(N4529), .A(a_man[19]), .B(N5163));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I942 (.Y(N5145), .A(N4896), .B(N4529));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1191 (.Y(N4274), .A0(N4634), .A1(N5115), .B0(N5145), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1472 (.Y(N4317), .A0(N4533), .A1(N13788), .B0(N4674), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1415 (.Y(N4924), .A0(N4533), .A1(N4314), .B0(N4341), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1519 (.Y(N5069), .A0(N4896), .A1(N4317), .B0(N4924), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1309 (.Y(N4734), .A0(N4533), .A1(N4849), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1355 (.Y(N4691), .A0(N4896), .A1(N4734), .B0(N4726), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1571 (.Y(N5156), .A0(N4634), .A1(N5069), .B0(N4691), .B1(a_man[21]));
AOI22X1 inst_cellmath__63_0_I5922 (.Y(N7339), .A0(a_man[22]), .A1(N4274), .B0(N4911), .B1(N5156));
INVX2 inst_cellmath__63_0_I1916 (.Y(N7533), .A(N7339));
NOR2XL inst_cellmath__63_0_I1955 (.Y(N7711), .A(N7350), .B(N7533));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1221 (.Y(N5010), .A0(N4314), .A1(N4869), .B0(N13752), .B1(N13786));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1463 (.Y(N5151), .A(N4533), .B(N5010));
INVXL inst_noninc_a_cellmath__55_2WWMM_I856 (.Y(N4582), .A(N4869));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1065 (.Y(N5064), .A0(N4479), .A1(N13807), .B0(N4736), .B1(N13786));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1406 (.Y(N4961), .A0(N4533), .A1(N4582), .B0(a_man[19]), .B1(N5064));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1510 (.Y(N5107), .A0(N4896), .A1(N5151), .B0(N4961), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1301 (.Y(N4771), .A0(N4533), .A1(N4154), .B0(N4519), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I868 (.Y(N4785), .A0(N13803), .A1(N4736), .B0(N4300), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1242 (.Y(N4442), .A0(N4533), .A1(N4785), .B0(N4489), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1346 (.Y(N4729), .A0(N4771), .A1(N4896), .B0(N4442), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1562 (.Y(N4171), .A0(N5107), .A1(N4634), .B0(N4729), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I866 (.Y(N4470), .A(N13806), .B(N4300));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I767 (.Y(N4390), .A0(N13797), .A1(N4953), .B0(N4300), .B1(N4826));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1083 (.Y(N4304), .A0(N4533), .A1(N4470), .B0(a_man[19]), .B1(N4390));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I991 (.Y(N4452), .A0(N13795), .A1(N13752), .B0(N4297), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1012 (.Y(N4242), .A0(N4533), .A1(N4452), .B0(a_man[19]), .B1(N4704));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1129 (.Y(N5150), .A0(N4896), .A1(N4304), .B0(a_man[20]), .B1(N4242));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I730 (.Y(N4402), .A(N4826), .B(N4438));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I886 (.Y(N4340), .A0(N5159), .A1(N4533), .B0(a_man[19]), .B1(N4402));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I787 (.Y(N4464), .A0(N4533), .A1(N4903), .B0(N4739), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I933 (.Y(N4164), .A0(N4896), .A1(N4340), .B0(N4464), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1182 (.Y(N4310), .A0(N4634), .A1(N5150), .B0(N4164), .B1(a_man[21]));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1614 (.Y(inst_cellmath__51[5]), .A0(N4911), .A1(N4171), .B0(a_man[22]), .B1(N4310));
INVX2 inst_cellmath__63_0_I1898 (.Y(N7627), .A(inst_cellmath__51[5]));
NOR2XL inst_cellmath__63_0_I2117 (.Y(N7086), .A(N3399), .B(N7627));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I727 (.Y(N4670), .A(N4826), .B(N4297));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1439 (.Y(N5075), .A0(N4314), .A1(N4438), .B0(N13760), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1466 (.Y(N5018), .A0(N4533), .A1(N4670), .B0(N5075), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1409 (.Y(N4607), .A0(N4470), .A1(N4533), .B0(a_man[19]), .B1(N5022));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1513 (.Y(N4750), .A0(N4896), .A1(N5018), .B0(N4607), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1274 (.Y(N4167), .A(N4314), .B(N4300));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1304 (.Y(N4420), .A0(N4167), .A1(N4533), .B0(a_man[19]), .B1(N4879));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1225 (.Y(N4741), .A(N4953), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1245 (.Y(N5113), .A0(N4741), .A1(N4533), .B0(a_man[19]), .B1(N13752));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1349 (.Y(N4375), .A0(N4896), .A1(N4420), .B0(N5113), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1565 (.Y(N4839), .A0(N4634), .A1(N4750), .B0(N4375), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1060 (.Y(N4822), .A0(N13806), .A1(N4297), .B0(a_man[17]), .B1(N13786));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1086 (.Y(N4966), .A(N4533), .B(N4822));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1015 (.Y(N4913), .A0(N4533), .A1(N4739), .B0(N4377), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1132 (.Y(N4796), .A0(N4966), .A1(N4896), .B0(a_man[20]), .B1(N4913));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I889 (.Y(N5002), .A0(N4533), .A1(N4390), .B0(a_man[19]), .B1(N4879));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I752 (.Y(N4190), .A0(N13795), .A1(N4953), .B0(N4736), .B1(N4826));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I722 (.Y(N5095), .A(N4314), .B(N4166));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I790 (.Y(N5137), .A0(N4533), .A1(N4190), .B0(N5095), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I936 (.Y(N4831), .A0(N4896), .A1(N5002), .B0(a_man[20]), .B1(N5137));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1185 (.Y(N4974), .A0(N4634), .A1(N4796), .B0(N4831), .B1(a_man[21]));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1617 (.Y(inst_cellmath__51[8]), .A0(N4911), .A1(N4839), .B0(N4974), .B1(a_man[22]));
INVX2 inst_cellmath__63_0_I1905 (.Y(N7594), .A(inst_cellmath__51[8]));
NOR2XL inst_cellmath__63_0_I2063 (.Y(N6997), .A(N3446), .B(N7594));
ADDFX1 inst_cellmath__63_0_I2318 (.CO(N6845), .S(N7536), .A(N7711), .B(N7086), .CI(N6997));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1383 (.Y(N4568), .A0(N4314), .A1(N4736), .B0(N4438), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I726 (.Y(N4981), .A0(N4314), .A1(N4479), .B0(a_man[17]), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1462 (.Y(N4931), .A0(N4533), .A1(N4568), .B0(N4981), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1384 (.Y(N5016), .A0(N4314), .A1(a_man[17]), .B0(N4869), .B1(N13782));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1405 (.Y(N4732), .A0(N4533), .A1(N5045), .B0(N5016), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1509 (.Y(N4882), .A0(N4931), .A1(N4896), .B0(a_man[20]), .B1(N4732));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1285 (.Y(N5121), .A0(N4314), .A1(N4869), .B0(N4300), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1300 (.Y(N4548), .A0(N4533), .A1(N5121), .B0(N4402), .B1(a_man[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I865 (.Y(N4598), .A(N13806), .B(N13745));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1241 (.Y(N4217), .A0(N4533), .A1(N4785), .B0(N4598), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1345 (.Y(N4509), .A0(N4548), .A1(N4896), .B0(N4217), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1561 (.Y(N4970), .A0(N4634), .A1(N4882), .B0(a_man[21]), .B1(N4509));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I979 (.Y(N4721), .A(N13795), .B(N4438));
AO22XL inst_noninc_a_cellmath__55_2WWMM_I871 (.Y(N4900), .A0(N13782), .A1(N4297), .B0(N13803), .B1(N4280));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I872 (.Y(N5127), .A(N4900));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1082 (.Y(N5099), .A0(N4721), .A1(N4533), .B0(a_man[19]), .B1(N5127));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1011 (.Y(N4595), .A(N4533), .B(N4489));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1128 (.Y(N4930), .A0(N4896), .A1(N5099), .B0(N4595), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I858 (.Y(N5026), .A(N4479), .B(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I885 (.Y(N5139), .A0(N5026), .A1(N4533), .B0(N4531), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I750 (.Y(N4325), .A0(N13795), .A1(N4736), .B0(N4953), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I716 (.Y(N4218), .A0(N4314), .A1(a_man[17]), .B0(N13745), .B1(N4826));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I786 (.Y(N4241), .A0(N4533), .A1(N4325), .B0(N4218), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I932 (.Y(N4962), .A0(N4896), .A1(N5139), .B0(N4241), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1181 (.Y(N5106), .A0(N4634), .A1(N4930), .B0(N4962), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1613 (.Y(inst_cellmath__51[4]), .A0(N4911), .A1(N4970), .B0(N5106), .B1(a_man[22]));
CLKBUFX2 inst_cellmath__63_0_I1894 (.Y(N6855), .A(inst_cellmath__51[4]));
INVX3 inst_cellmath__63_0_I1895 (.Y(N7050), .A(N6855));
NOR2XL inst_cellmath__63_0_I2135 (.Y(N7117), .A(N3432), .B(N7050));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1467 (.Y(N4221), .A0(N4533), .A1(N4939), .B0(N4929), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1061 (.Y(N4250), .A0(N13763), .A1(N13806), .B0(N13786), .B1(N13745));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1410 (.Y(N4830), .A0(N4533), .A1(N4250), .B0(N4822), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1514 (.Y(N4975), .A0(N4896), .A1(N4221), .B0(a_man[20]), .B1(N4830));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I831 (.Y(N4308), .A0(N13797), .A1(N4280), .B0(N13754), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1305 (.Y(N4647), .A0(N4533), .A1(N5163), .B0(N4308), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1246 (.Y(N4316), .A0(N4533), .A1(N4875), .B0(N5081), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1350 (.Y(N4602), .A0(N4896), .A1(N4647), .B0(N4316), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1566 (.Y(N5063), .A0(N4634), .A1(N4975), .B0(N4602), .B1(a_man[21]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1087 (.Y(N4391), .A(a_man[19]), .B(N4469));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1016 (.Y(N5138), .A0(N4768), .A1(N4533), .B0(a_man[19]), .B1(N5045));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1133 (.Y(N5017), .A0(N4896), .A1(N4391), .B0(N5138), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I890 (.Y(N4205), .A0(N4533), .A1(N4540), .B0(N4308), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I753 (.Y(N4411), .A0(N13791), .A1(N4280), .B0(N4438), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I791 (.Y(N4337), .A0(N4533), .A1(N4411), .B0(N13745), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I937 (.Y(N5053), .A0(N4896), .A1(N4205), .B0(N4337), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1186 (.Y(N4175), .A0(N4634), .A1(N5017), .B0(N5053), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1618 (.Y(inst_cellmath__51[9]), .A0(N4911), .A1(N5063), .B0(N4175), .B1(a_man[22]));
INVX2 inst_cellmath__63_0_I1907 (.Y(N7288), .A(inst_cellmath__51[9]));
NOR2XL inst_cellmath__63_0_I2045 (.Y(N6966), .A(N3412), .B(N7288));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I970 (.Y(N4599), .A0(N4280), .A1(N13803), .B0(N13772), .B1(N13745));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1468 (.Y(N4444), .A0(N4533), .A1(N4741), .B0(N4599), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1411 (.Y(N5051), .A0(N4533), .A1(N4540), .B0(N4469), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1515 (.Y(N4176), .A0(N4444), .A1(N4896), .B0(a_man[20]), .B1(N5051));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1306 (.Y(N4868), .A0(N4533), .A1(N4413), .B0(N5124), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1247 (.Y(N4530), .A0(N4533), .A1(N5081), .B0(N5127), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1351 (.Y(N4823), .A0(N4896), .A1(N4868), .B0(N4530), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1567 (.Y(N4269), .A0(N4634), .A1(N4176), .B0(N4823), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1088 (.Y(N5059), .A0(N4533), .A1(N4250), .B0(N13752), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1017 (.Y(N4338), .A0(N4533), .A1(N4805), .B0(N4471), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1134 (.Y(N4220), .A0(N4896), .A1(N5059), .B0(a_man[20]), .B1(N4338));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I863 (.Y(N4988), .A0(N13806), .A1(N4300), .B0(N4438), .B1(N13782));
INVX1 inst_noninc_a_cellmath__55_2WWMM_I5799 (.Y(N13764), .A(N13761));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I832 (.Y(N4747), .A0(N13806), .A1(N13764), .B0(a_man[17]), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I891 (.Y(N4424), .A0(N4988), .A1(N4533), .B0(a_man[19]), .B1(N4747));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I792 (.Y(N4549), .A0(N4533), .A1(N5081), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I938 (.Y(N4257), .A0(N4896), .A1(N4424), .B0(N4549), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1187 (.Y(N4396), .A0(N4634), .A1(N4220), .B0(N4257), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1619 (.Y(inst_cellmath__51[10]), .A0(N4911), .A1(N4269), .B0(N4396), .B1(a_man[22]));
INVX2 inst_cellmath__63_0_I1909 (.Y(N6983), .A(inst_cellmath__51[10]));
NOR2XL inst_cellmath__63_0_I2027 (.Y(N6940), .A(N3456), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2321 (.CO(N7118), .S(N6921), .A(N7117), .B(N6966), .CI(N6940));
ADDFX1 inst_cellmath__63_0_I2337 (.CO(N7098), .S(N6903), .A(N7614), .B(N6845), .CI(N7118));
ADDFX1 inst_cellmath__63_0_I2325 (.CO(N6889), .S(N7580), .A(N7421), .B(N7536), .CI(N6921));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1473 (.Y(N4532), .A(N4644), .B(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1520 (.Y(N4275), .A0(N4896), .A1(N4532), .B0(N4718), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1356 (.Y(N4920), .A0(N4896), .A1(N4934), .B0(N4726), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1572 (.Y(N4356), .A0(N4634), .A1(N4275), .B0(N4920), .B1(a_man[21]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1192 (.Y(N4926), .A(N4896), .B(N4692));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1193 (.Y(N4494), .A(N4926), .B(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1624 (.Y(inst_cellmath__51[15]), .A0(N4911), .A1(N4356), .B0(N4494), .B1(a_man[22]));
INVX2 inst_cellmath__63_0_I1918 (.Y(N7304), .A(inst_cellmath__51[15]));
NOR2XL inst_cellmath__63_0_I1956 (.Y(N7206), .A(N7350), .B(N7304));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I749 (.Y(N5122), .A0(N13795), .A1(N4166), .B0(N4826), .B1(N4953));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1460 (.Y(N4485), .A0(N4533), .A1(N5122), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1403 (.Y(N4295), .A0(N4533), .A1(N4582), .B0(N4568), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1507 (.Y(N4434), .A0(N4896), .A1(N4485), .B0(a_man[20]), .B1(N4295));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1283 (.Y(N4227), .A0(N4438), .A1(N4314), .B0(N4280), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1272 (.Y(N4949), .A0(N4314), .A1(N4438), .B0(N13745), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1298 (.Y(N5136), .A0(N4227), .A1(N4533), .B0(a_man[19]), .B1(N4949));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I715 (.Y(N4794), .A0(N4314), .A1(N4300), .B0(N4736), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1239 (.Y(N4793), .A0(N4533), .A1(N4794), .B0(a_man[19]), .B1(N4747));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1343 (.Y(N5085), .A0(N4896), .A1(N5136), .B0(N4793), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1559 (.Y(N4521), .A0(N4634), .A1(N4434), .B0(a_man[21]), .B1(N5085));
INVXL inst_noninc_a_cellmath__55_2WWMM_I1049 (.Y(N4520), .A(N4280));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1080 (.Y(N4654), .A0(N4533), .A1(N4721), .B0(N4520), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I989 (.Y(N4802), .A0(N13795), .A1(N13763), .B0(N4438), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1009 (.Y(N4150), .A0(N4533), .A1(N4802), .B0(a_man[19]), .B1(N4599));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1126 (.Y(N4484), .A0(N4896), .A1(N4654), .B0(a_man[20]), .B1(N4150));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I825 (.Y(N4743), .A0(N13797), .A1(N4166), .B0(N4280), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I883 (.Y(N4689), .A0(N4582), .A1(N4533), .B0(N4743), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I748 (.Y(N4894), .A0(N13795), .A1(N13762), .B0(N4826), .B1(N4166));
INVXL inst_noninc_a_cellmath__55_2WWMM_I714 (.Y(N4779), .A(N4300));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I784 (.Y(N4815), .A0(N4533), .A1(N4894), .B0(N4779), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I930 (.Y(N4513), .A0(N4896), .A1(N4689), .B0(N4815), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1179 (.Y(N4659), .A0(N4634), .A1(N4484), .B0(N4513), .B1(a_man[21]));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1611 (.Y(inst_cellmath__51[2]), .A0(N4911), .A1(N4521), .B0(a_man[22]), .B1(N4659));
INVX2 inst_cellmath__63_0_I1890 (.Y(N7663), .A(inst_cellmath__51[2]));
NOR2XL inst_cellmath__63_0_I2190 (.Y(N7585), .A(N3538), .B(N7663));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1464 (.Y(N4570), .A0(N4533), .A1(N4496), .B0(a_man[17]), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1288 (.Y(N4170), .A0(N4314), .A1(N4300), .B0(N4869), .B1(N13782));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1407 (.Y(N4163), .A0(N4533), .A1(N4177), .B0(N4170), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1511 (.Y(N4311), .A0(N4896), .A1(N4570), .B0(a_man[20]), .B1(N4163));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1000 (.Y(N4969), .A0(N13752), .A1(N13806), .B0(N13763), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I869 (.Y(N4428), .A0(N4280), .A1(N13803), .B0(N4166), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1302 (.Y(N4996), .A0(N4533), .A1(N4969), .B0(N4428), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1223 (.Y(N4652), .A(N13760), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1218 (.Y(N4592), .A0(N13803), .A1(N13752), .B0(a_man[17]), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1243 (.Y(N4665), .A0(N4533), .A1(N4652), .B0(N4592), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1347 (.Y(N4956), .A0(N4896), .A1(N4996), .B0(N4665), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1563 (.Y(N4393), .A0(N4634), .A1(N4311), .B0(N4956), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1084 (.Y(N4518), .A0(N4533), .A1(N4517), .B0(a_man[19]), .B1(N4392));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I974 (.Y(N4354), .A0(N13752), .A1(N13791), .B0(N13772), .B1(N4869));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1013 (.Y(N4466), .A0(N4271), .A1(N4533), .B0(N4354), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1130 (.Y(N4351), .A0(N4896), .A1(N4518), .B0(a_man[20]), .B1(N4466));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I827 (.Y(N5060), .A(N4826), .B(N4479));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I887 (.Y(N4554), .A0(N4533), .A1(N4897), .B0(N5060), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I717 (.Y(N4650), .A0(N4314), .A1(N4995), .B0(N4736), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I788 (.Y(N4686), .A0(N4533), .A1(N4218), .B0(N4650), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I934 (.Y(N4383), .A0(N4896), .A1(N4554), .B0(N4686), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1183 (.Y(N4524), .A0(N4634), .A1(N4351), .B0(N4383), .B1(a_man[21]));
AOI22X2 inst_noninc_a_cellmath__55_2WWMM_I1615 (.Y(inst_cellmath__51[6]), .A0(N4911), .A1(N4393), .B0(N4524), .B1(a_man[22]));
INVX3 inst_cellmath__63_0_I1900 (.Y(N7321), .A(inst_cellmath__51[6]));
NOR2XL inst_cellmath__63_0_I2118 (.Y(N7473), .A(N3399), .B(N7321));
ADDFX1 inst_cellmath__63_0_I2333 (.CO(N7320), .S(N7129), .A(N7206), .B(N7585), .CI(N7473));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1438 (.Y(N4226), .A(N4166), .B(N13782));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1459 (.Y(N4263), .A0(N4533), .A1(N4162), .B0(N4226), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I820 (.Y(N4561), .A0(N13803), .A1(N4869), .B0(N4297), .B1(N4826));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1402 (.Y(N5089), .A0(N4533), .A1(N4457), .B0(N4561), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1506 (.Y(N4213), .A0(N4896), .A1(N4263), .B0(N5089), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1282 (.Y(N5024), .A0(N4314), .A1(N13745), .B0(N13760), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1297 (.Y(N4909), .A0(N4533), .A1(N5024), .B0(N4344), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I995 (.Y(N4557), .A0(N13807), .A1(N4479), .B0(N4280), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I854 (.Y(N5158), .A0(N4736), .A1(N13803), .B0(N13782), .B1(N4166));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1238 (.Y(N4566), .A0(N4533), .A1(N4557), .B0(N5158), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1342 (.Y(N4861), .A0(N4896), .A1(N4909), .B0(N4566), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1558 (.Y(N4305), .A0(N4634), .A1(N4213), .B0(N4861), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1059 (.Y(N4194), .A0(N13806), .A1(N4479), .B0(N4297), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1079 (.Y(N4427), .A0(N4533), .A1(N4194), .B0(N4471), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I733 (.Y(N4717), .A0(N4314), .A1(N4736), .B0(N4869), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1008 (.Y(N4950), .A0(N4533), .A1(N4717), .B0(N5127), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1125 (.Y(N4262), .A0(N4896), .A1(N4427), .B0(N4950), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I882 (.Y(N4467), .A0(N4533), .A1(N4674), .B0(N4162), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I747 (.Y(N4450), .A(N13795), .B(N13744));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I713 (.Y(N4553), .A0(N4314), .A1(N13760), .B0(N13745), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I783 (.Y(N4593), .A0(N4533), .A1(N4450), .B0(N4553), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I929 (.Y(N4296), .A0(N4896), .A1(N4467), .B0(N4593), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1178 (.Y(N4433), .A0(N4634), .A1(N4262), .B0(N4296), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1610 (.Y(inst_cellmath__51[1]), .A0(N4911), .A1(N4305), .B0(N4433), .B1(a_man[22]));
NAND2XL inst_cellmath__63_0_I2208 (.Y(N7615), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[1]));
INVXL inst_cellmath__63_0_I1921 (.Y(N6885), .A(a_man[0]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1521 (.Y(N4495), .A(N4896), .B(N5074));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1357 (.Y(N5143), .A(N4726), .B(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1573 (.Y(N4580), .A0(N4634), .A1(N4495), .B0(N5143), .B1(a_man[21]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1625 (.Y(inst_cellmath__51[16]), .A(a_man[22]), .B(N4580));
INVXL inst_cellmath__63_0_I1919 (.Y(N6998), .A(inst_cellmath__51[16]));
NOR2XL inst_cellmath__63_0_I1938 (.Y(N7180), .A(N6885), .B(N6998));
NOR2XL inst_cellmath__63_0_I2100 (.Y(N7442), .A(N3702), .B(N7016));
ADDFX1 inst_cellmath__63_0_I2331 (.CO(N7433), .S(N7237), .A(N7615), .B(N7180), .CI(N7442));
NOR2XL inst_cellmath__63_0_I1992 (.Y(N7264), .A(N3603), .B(N6952));
NOR2XL inst_cellmath__63_0_I1974 (.Y(N7235), .A(N3142), .B(N7533));
NOR2XL inst_cellmath__63_0_I2010 (.Y(N7296), .A(N7257), .B(N3503));
ADDFXL inst_cellmath__63_0_I2334 (.CO(N7708), .S(N7517), .A(N7264), .B(N7235), .CI(N7296));
ADDFXL inst_cellmath__63_0_I2338 (.CO(N7485), .S(N7287), .A(N7129), .B(N7237), .CI(N7517));
ADDFXL inst_cellmath__63_0_I2341 (.CO(N6870), .S(N7561), .A(N6903), .B(N6889), .CI(N7287));
NOR2XL inst_cellmath__63_0_I1936 (.Y(N7292), .A(N6885), .B(N7533));
NOR2XL inst_cellmath__63_0_I2152 (.Y(N7643), .A(N3462), .B(N7663));
NOR2XL inst_cellmath__63_0_I1954 (.Y(N7323), .A(N7350), .B(N6952));
ADDFX1 inst_cellmath__63_0_I2304 (.CO(N7631), .S(N7439), .A(N7292), .B(N7643), .CI(N7323));
INVXL inst_noninc_a_cellmath__55_2WWMM_I1446 (.Y(N4371), .A(N4479));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I985 (.Y(N4998), .A0(N4280), .A1(N13795), .B0(N4479), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1458 (.Y(N5057), .A0(N4533), .A1(N4371), .B0(N4998), .B1(a_man[19]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I1382 (.Y(N5149), .A(N4736));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1401 (.Y(N4865), .A0(N4533), .A1(N5158), .B0(N5149), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1505 (.Y(N5009), .A0(N4896), .A1(N5057), .B0(N4865), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1281 (.Y(N4579), .A(N4314), .B(N4297));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1271 (.Y(N4286), .A(N13745), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1296 (.Y(N4685), .A0(N4533), .A1(N4579), .B0(N4286), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I723 (.Y(N4572), .A0(N4314), .A1(N4995), .B0(N4300), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1237 (.Y(N4348), .A0(N4533), .A1(N4572), .B0(N4786), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1341 (.Y(N4642), .A0(N4896), .A1(N4685), .B0(N4348), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1557 (.Y(N5103), .A0(N4634), .A1(N5009), .B0(N4642), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1048 (.Y(N5102), .A0(N13795), .A1(N4736), .B0(N13745), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1078 (.Y(N4208), .A0(N4533), .A1(N4802), .B0(N5102), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I969 (.Y(N4616), .A0(N13803), .A1(N4736), .B0(N4297), .B1(N13772));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1007 (.Y(N4723), .A0(N4533), .A1(N4252), .B0(N4616), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1124 (.Y(N5056), .A0(N4208), .A1(N4896), .B0(a_man[20]), .B1(N4723));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I881 (.Y(N4244), .A0(N4533), .A1(N5158), .B0(N4561), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I712 (.Y(N4339), .A0(N4314), .A1(N4736), .B0(a_man[17]), .B1(N4826));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I782 (.Y(N4366), .A0(N4533), .A1(N4457), .B0(a_man[19]), .B1(N4339));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I928 (.Y(N5090), .A0(N4896), .A1(N4244), .B0(a_man[20]), .B1(N4366));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1177 (.Y(N4212), .A0(N4634), .A1(N5056), .B0(N5090), .B1(a_man[21]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1609 (.Y(inst_cellmath__51[0]), .A0(N5103), .A1(N4911), .B0(a_man[22]), .B1(N4212));
NAND2XL inst_cellmath__63_0_I2207 (.Y(N7226), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[0]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1440 (.Y(N4550), .A0(N4314), .A1(N4280), .B0(N4869), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1461 (.Y(N4701), .A0(N4533), .A1(N4550), .B0(N4286), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1389 (.Y(N4243), .A0(N4314), .A1(N4438), .B0(N4479), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1404 (.Y(N4512), .A0(N4533), .A1(N4243), .B0(N4584), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1508 (.Y(N4660), .A0(N4896), .A1(N4701), .B0(N4512), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1284 (.Y(N4449), .A(N4314), .B(N13766));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I988 (.Y(N4656), .A0(N13795), .A1(N13764), .B0(N13782), .B1(N4297));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1299 (.Y(N4336), .A0(N4533), .A1(N4449), .B0(N4656), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1240 (.Y(N5014), .A0(N4533), .A1(N4354), .B0(N4875), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1344 (.Y(N4293), .A0(N4896), .A1(N4336), .B0(N5014), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1560 (.Y(N4744), .A0(N4634), .A1(N4660), .B0(N4293), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1081 (.Y(N4876), .A0(N4354), .A1(N4533), .B0(a_man[19]), .B1(N4615));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I971 (.Y(N4266), .A0(N13752), .A1(N13803), .B0(N13772), .B1(N4736));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1010 (.Y(N4368), .A0(N4533), .A1(N5101), .B0(a_man[19]), .B1(N4266));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1127 (.Y(N4700), .A0(N4896), .A1(N4876), .B0(a_man[20]), .B1(N4368));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I857 (.Y(N4804), .A0(N13806), .A1(N4438), .B0(N4736), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I826 (.Y(N4967), .A0(N13797), .A1(N4479), .B0(N13745), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I884 (.Y(N4914), .A0(N4804), .A1(N4533), .B0(a_man[19]), .B1(N4967));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I785 (.Y(N5039), .A0(N4533), .A1(N5122), .B0(a_man[19]), .B1(N4794));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I931 (.Y(N4733), .A0(N4896), .A1(N4914), .B0(N5039), .B1(a_man[20]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1180 (.Y(N4881), .A0(N4634), .A1(N4700), .B0(N4733), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1612 (.Y(inst_cellmath__51[3]), .A0(N4911), .A1(N4744), .B0(a_man[22]), .B1(N4881));
CLKBUFX2 inst_cellmath__63_0_I1892 (.Y(N7159), .A(inst_cellmath__51[3]));
INVX3 inst_cellmath__63_0_I1893 (.Y(N7354), .A(N7159));
NOR2XL inst_cellmath__63_0_I2153 (.Y(N7146), .A(N3462), .B(N7354));
XNOR2X1 inst_cellmath__63_0_I2316 (.Y(N7647), .A(N7226), .B(N7146));
NOR2XL inst_cellmath__63_0_I2080 (.Y(N7527), .A(N3611), .B(N7321));
NOR2XL inst_cellmath__63_0_I2044 (.Y(N7470), .A(N3412), .B(N7594));
NOR2XL inst_cellmath__63_0_I2116 (.Y(N7583), .A(N3399), .B(N7050));
ADDFX1 inst_cellmath__63_0_I2306 (.CO(N7522), .S(N7326), .A(N7527), .B(N7470), .CI(N7583));
ADDFX1 inst_cellmath__63_0_I2323 (.CO(N7002), .S(N7695), .A(N7631), .B(N7647), .CI(N7522));
INVX1 inst_cellmath__63_0_I1886 (.Y(N7085), .A(inst_cellmath__51[1]));
NOR2XL inst_cellmath__63_0_I2151 (.Y(N7255), .A(N3462), .B(N7085));
INVX1 inst_cellmath__63_0_I1884 (.Y(N7310), .A(inst_cellmath__51[0]));
NOR2XL inst_cellmath__63_0_I2169 (.Y(N7282), .A(N3496), .B(N7310));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1469 (.Y(N4668), .A0(N4533), .A1(N5095), .B0(N13760), .B1(a_man[19]));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1412 (.Y(N4256), .A0(N4457), .A1(N4533), .B0(a_man[19]), .B1(N4268));
AOI22X1 inst_noninc_a_cellmath__55_2WWMM_I1516 (.Y(N4397), .A0(N4668), .A1(N4896), .B0(a_man[20]), .B1(N4256));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1307 (.Y(N5091), .A0(N4533), .A1(N13745), .B0(N4802), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1248 (.Y(N4755), .A0(N4533), .A1(N4988), .B0(N5022), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1352 (.Y(N5047), .A0(N4896), .A1(N5091), .B0(N4755), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1568 (.Y(N4491), .A0(N4634), .A1(N4397), .B0(N5047), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1089 (.Y(N4267), .A0(N4533), .A1(N4540), .B0(N5081), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I766 (.Y(N4958), .A0(a_man[17]), .A1(N13797), .B0(N13762), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1018 (.Y(N4552), .A0(N4533), .A1(N5045), .B0(N4958), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1135 (.Y(N4443), .A0(N4896), .A1(N4267), .B0(N4552), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I794 (.Y(N4772), .A0(N4533), .A1(N4768), .B0(N13788), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I939 (.Y(N4478), .A0(N4896), .A1(N4651), .B0(N4772), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1188 (.Y(N4621), .A0(N4634), .A1(N4443), .B0(N4478), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1620 (.Y(inst_cellmath__51[11]), .A0(N4911), .A1(N4491), .B0(N4621), .B1(a_man[22]));
INVX1 inst_cellmath__63_0_I1910 (.Y(N7562), .A(inst_cellmath__51[11]));
NOR2XL inst_cellmath__63_0_I1971 (.Y(N6963), .A(N3142), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2295 (.CO(N7698), .S(N7508), .A(N7255), .B(N7282), .CI(N6963));
ADDFX1 inst_cellmath__63_0_I2310 (.CO(N7291), .S(N7102), .A(N7439), .B(N7698), .CI(N7326));
NOR2XL inst_cellmath__63_0_I2188 (.Y(N7699), .A(N3538), .B(N7310));
NOR2XL inst_cellmath__63_0_I2008 (.Y(N7409), .A(N3503), .B(N6983));
NOR2X1 inst_cellmath__63_0_I2170 (.Y(N7673), .A(N3496), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2307 (.CO(N7020), .S(N6832), .A(N7699), .B(N7409), .CI(N7673));
NOR2XL inst_cellmath__63_0_I2062 (.Y(N7500), .A(N3446), .B(N7016));
NOR2XL inst_cellmath__63_0_I2134 (.Y(N7613), .A(N3432), .B(N7354));
NOR2XL inst_cellmath__63_0_I2026 (.Y(N7440), .A(N3456), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2305 (.CO(N7135), .S(N6939), .A(N7500), .B(N7613), .CI(N7440));
NOR2XL inst_cellmath__63_0_I2171 (.Y(N7170), .A(N3496), .B(N7663));
NOR2XL inst_cellmath__63_0_I1937 (.Y(N7681), .A(N6885), .B(N7304));
NOR2X1 inst_cellmath__63_0_I2099 (.Y(N7058), .A(N3702), .B(N7321));
ADDFXL inst_cellmath__63_0_I2319 (.CO(N7225), .S(N7036), .A(N7681), .B(N7058), .CI(N7170));
ADDFX1 inst_cellmath__63_0_I2324 (.CO(N7385), .S(N7193), .A(N7020), .B(N7135), .CI(N7036));
ADDFX1 inst_cellmath__63_0_I2327 (.CO(N7662), .S(N7469), .A(N7695), .B(N7291), .CI(N7193));
NOR2XL inst_cellmath__63_0_I2079 (.Y(N7143), .A(N3611), .B(N7627));
NOR2XL inst_cellmath__63_0_I1953 (.Y(N6936), .A(N7350), .B(N7257));
ADDHX1 inst_cellmath__63_0_I2291 (.CO(N7040), .S(N6846), .A(N7143), .B(N6936));
NOR2XL inst_cellmath__63_0_I2060 (.Y(N7611), .A(N3446), .B(N7627));
NOR2XL inst_cellmath__63_0_I1934 (.Y(N7406), .A(N6885), .B(N7257));
ADDHX1 inst_cellmath__63_0_I2280 (.CO(N7215), .S(N7025), .A(N7611), .B(N7406));
NOR2XL inst_cellmath__63_0_I2006 (.Y(N7526), .A(N3503), .B(N7594));
NOR2XL inst_cellmath__63_0_I2024 (.Y(N7550), .A(N3456), .B(N7016));
NOR2XL inst_cellmath__63_0_I1970 (.Y(N7467), .A(N3142), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2282 (.CO(N7106), .S(N6911), .A(N7526), .B(N7550), .CI(N7467));
ADDFXL inst_cellmath__63_0_I2296 (.CO(N7198), .S(N7006), .A(N6846), .B(N7215), .CI(N7106));
ADDFX1 inst_cellmath__63_0_I2311 (.CO(N7679), .S(N7488), .A(N6832), .B(N6939), .CI(N7198));
NOR2XL inst_cellmath__63_0_I2078 (.Y(N7640), .A(N3611), .B(N7050));
NOR2XL inst_cellmath__63_0_I2042 (.Y(N7581), .A(N3412), .B(N7321));
NOR2XL inst_cellmath__63_0_I2150 (.Y(N6869), .A(N3462), .B(N7310));
ADDFX1 inst_cellmath__63_0_I2283 (.CO(N7491), .S(N7295), .A(N7640), .B(N7581), .CI(N6869));
NOR2XL inst_cellmath__63_0_I2096 (.Y(N7670), .A(N3702), .B(N7354));
NOR2XL inst_cellmath__63_0_I2114 (.Y(N7696), .A(N3399), .B(N7663));
NOR2XL inst_cellmath__63_0_I1988 (.Y(N7495), .A(N3603), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2281 (.CO(N7603), .S(N7408), .A(N7670), .B(N7696), .CI(N7495));
NOR2X1 inst_cellmath__63_0_I2115 (.Y(N7197), .A(N7354), .B(N3399));
NOR2XL inst_cellmath__63_0_I2133 (.Y(N7224), .A(N3432), .B(N7663));
NOR2XL inst_cellmath__63_0_I2007 (.Y(N7026), .A(N3503), .B(N7288));
ADDFXL inst_cellmath__63_0_I2292 (.CO(N7423), .S(N7228), .A(N7224), .B(N7197), .CI(N7026));
ADDFXL inst_cellmath__63_0_I2297 (.CO(N7584), .S(N7389), .A(N7491), .B(N7603), .CI(N7228));
NOR2XL inst_cellmath__63_0_I1990 (.Y(N7379), .A(N3603), .B(N7562));
NOR2XL inst_cellmath__63_0_I2098 (.Y(N7551), .A(N3702), .B(N7627));
NOR2XL inst_cellmath__63_0_I1972 (.Y(N7349), .A(N3142), .B(N7257));
ADDHX1 inst_cellmath__63_0_I2303 (.CO(N7243), .S(N7055), .A(N7551), .B(N7349));
ADDFX1 inst_cellmath__63_0_I2308 (.CO(N7404), .S(N7210), .A(N7040), .B(N7379), .CI(N7055));
NOR2XL inst_cellmath__63_0_I2097 (.Y(N7167), .A(N3702), .B(N7050));
NOR2XL inst_cellmath__63_0_I2061 (.Y(N7114), .A(N3446), .B(N7321));
NOR2XL inst_cellmath__63_0_I1935 (.Y(N6909), .A(N6885), .B(N6952));
ADDFXL inst_cellmath__63_0_I2294 (.CO(N7313), .S(N7122), .A(N7167), .B(N7114), .CI(N6909));
NOR2XL inst_cellmath__63_0_I2025 (.Y(N7056), .A(N3456), .B(N7594));
NOR2XL inst_cellmath__63_0_I2043 (.Y(N7083), .A(N3412), .B(N7016));
NOR2XL inst_cellmath__63_0_I1989 (.Y(N6995), .A(N3603), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2293 (.CO(N6925), .S(N7617), .A(N7056), .B(N7083), .CI(N6995));
NOR2XL inst_cellmath__63_0_I2132 (.Y(N6844), .A(N3432), .B(N7085));
NOR2XL inst_cellmath__63_0_I1952 (.Y(N7436), .A(N7350), .B(N7562));
NOR2XL inst_cellmath__63_0_I2041 (.Y(N7194), .A(N3412), .B(N7627));
NOR2XL inst_cellmath__63_0_I1951 (.Y(N7052), .A(N7350), .B(N6983));
ADDHX1 inst_cellmath__63_0_I2270 (.CO(N6899), .S(N7588), .A(N7194), .B(N7052));
ADDFX1 inst_cellmath__63_0_I2284 (.CO(N6989), .S(N7683), .A(N6844), .B(N7436), .CI(N6899));
ADDFX1 inst_cellmath__63_0_I2298 (.CO(N7088), .S(N6894), .A(N7122), .B(N7617), .CI(N6989));
ADDFXL inst_cellmath__63_0_I2312 (.CO(N7178), .S(N6985), .A(N7584), .B(N7210), .CI(N7088));
ADDFX1 inst_cellmath__63_0_I2328 (.CO(N7158), .S(N6965), .A(N7580), .B(N7679), .CI(N7178));
ADDFX1 inst_cellmath__63_0_I2343 (.CO(N7644), .S(N7452), .A(N7561), .B(N7662), .CI(N7158));
OR2XL inst_cellmath__63_0_I2317 (.Y(N6954), .A(N7226), .B(N7146));
NOR2XL inst_cellmath__63_0_I2028 (.Y(N7327), .A(N3456), .B(N7562));
ADDFXL inst_cellmath__63_0_I2336 (.CO(N7593), .S(N7398), .A(N6954), .B(N7327), .CI(N7225));
ADDFXL inst_cellmath__63_0_I2340 (.CO(N7369), .S(N7175), .A(N7398), .B(N7002), .CI(N7385));
NOR2XL inst_cellmath__63_0_I2173 (.Y(N7061), .A(N3496), .B(N7050));
NOR2XL inst_cellmath__63_0_I2011 (.Y(N7684), .A(N3503), .B(N6952));
NOR2XL inst_cellmath__63_0_I2029 (.Y(N6833), .A(N3456), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2349 (.CO(N7303), .S(N7113), .A(N7061), .B(N7684), .CI(N6833));
NOR2XL inst_cellmath__63_0_I2119 (.Y(N6969), .A(N3399), .B(N7016));
NOR2XL inst_cellmath__63_0_I1993 (.Y(N7655), .A(N3603), .B(N7533));
NOR2XL inst_cellmath__63_0_I2083 (.Y(N6914), .A(N3611), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2347 (.CO(N7416), .S(N7221), .A(N6969), .B(N7655), .CI(N6914));
ADDFX1 inst_cellmath__63_0_I2353 (.CO(N7079), .S(N6883), .A(N7113), .B(N7221), .CI(N7593));
ADDFXL inst_cellmath__63_0_I2356 (.CO(N7348), .S(N7155), .A(N7369), .B(N6883), .CI(N6870));
NAND2XL inst_cellmath__63_0_I2209 (.Y(N7120), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[2]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1358 (.Y(N4560), .A(N4896), .B(N4529));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I1626 (.Y(inst_cellmath__51[17]), .A0N(N4560), .A1N(a_man[21]), .B0(N4911));
INVXL inst_cellmath__63_0_I1920 (.Y(N7576), .A(inst_cellmath__51[17]));
NOR2XL inst_cellmath__63_0_I1939 (.Y(N7565), .A(N6885), .B(N7576));
NOR2XL inst_cellmath__63_0_I1957 (.Y(N7596), .A(N7350), .B(N6998));
ADDFX1 inst_cellmath__63_0_I2345 (.CO(N7532), .S(N7337), .A(N7565), .B(N7596), .CI(N7120));
ADDFX1 inst_cellmath__63_0_I2351 (.CO(N7190), .S(N6996), .A(N7320), .B(N7337), .CI(N7708));
NOR2XL inst_cellmath__63_0_I2154 (.Y(N7531), .A(N3462), .B(N7050));
NOR2XL inst_cellmath__63_0_I2064 (.Y(N7382), .A(N3446), .B(N7288));
NOR2XL inst_cellmath__63_0_I2046 (.Y(N7352), .A(N3412), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2335 (.CO(N7204), .S(N7015), .A(N7382), .B(N7531), .CI(N7352));
NOR2XL inst_cellmath__63_0_I2172 (.Y(N7555), .A(N7354), .B(N3496));
NOR2XL inst_cellmath__63_0_I2136 (.Y(N7503), .A(N3432), .B(N7627));
NOR2XL inst_cellmath__63_0_I2082 (.Y(N7411), .A(N3611), .B(N7594));
ADDFX1 inst_cellmath__63_0_I2332 (.CO(N6934), .S(N7626), .A(N7555), .B(N7503), .CI(N7411));
NOR2XL inst_cellmath__63_0_I2189 (.Y(N7199), .A(N3538), .B(N7085));
NOR2XL inst_cellmath__63_0_I2009 (.Y(N6912), .A(N3503), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2322 (.CO(N7504), .S(N7308), .A(N7199), .B(N6912), .CI(N7243));
ADDFX1 inst_cellmath__63_0_I2339 (.CO(N6982), .S(N7677), .A(N7015), .B(N7626), .CI(N7504));
NOR2XL inst_cellmath__63_0_I1975 (.Y(N7622), .A(N3142), .B(N7304));
NOR2XL inst_cellmath__63_0_I2155 (.Y(N7031), .A(N3462), .B(N7627));
NOR2X1 inst_cellmath__63_0_I2137 (.Y(N7001), .A(N3432), .B(N7321));
ADDFX1 inst_cellmath__63_0_I2346 (.CO(N7032), .S(N6841), .A(N7001), .B(N7622), .CI(N7031));
NOR2X1 inst_cellmath__63_0_I2191 (.Y(N7090), .A(N3538), .B(N7354));
NOR2XL inst_cellmath__63_0_I2101 (.Y(N6941), .A(N3702), .B(N7594));
NOR2XL inst_cellmath__63_0_I2065 (.Y(N6884), .A(N3446), .B(N6983));
ADDFXL inst_cellmath__63_0_I2348 (.CO(N6919), .S(N7610), .A(N7090), .B(N6941), .CI(N6884));
ADDFXL inst_cellmath__63_0_I2352 (.CO(N7575), .S(N7381), .A(N6841), .B(N7204), .CI(N7610));
ADDFXL inst_cellmath__63_0_I2355 (.CO(N6962), .S(N7657), .A(N6996), .B(N6982), .CI(N7381));
NOR2XL inst_cellmath__63_0_I2047 (.Y(N6854), .A(N3412), .B(N7562));
ADDFXL inst_cellmath__63_0_I2350 (.CO(N7691), .S(N7499), .A(N7433), .B(N6854), .CI(N6934));
ADDFX1 inst_cellmath__63_0_I2354 (.CO(N7465), .S(N7265), .A(N7499), .B(N7098), .CI(N7485));
ADDFX1 inst_cellmath__63_0_I2309 (.CO(N6907), .S(N7599), .A(N6925), .B(N7423), .CI(N7313));
ADDFX1 inst_cellmath__63_0_I2326 (.CO(N7270), .S(N7084), .A(N7308), .B(N7404), .CI(N6907));
ADDFXL inst_cellmath__63_0_I2342 (.CO(N7256), .S(N7066), .A(N7677), .B(N7270), .CI(N7175));
ADDFXL inst_cellmath__63_0_I2357 (.CO(N6850), .S(N7541), .A(N7657), .B(N7265), .CI(N7256));
ADDFXL inst_cellmath__64_0_I16112 (.CO(inst_cellmath__63__W0[18]), .S(N26263), .A(N7644), .B(N7155), .CI(N7541));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1219 (.Y(N4382), .A0(N4314), .A1(N4953), .B0(N4297), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1441 (.Y(N4773), .A0(N4314), .A1(N4300), .B0(N13754), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1477 (.Y(N5073), .A0(N4533), .A1(N4382), .B0(N4773), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1386 (.Y(N4363), .A0(N4314), .A1(N13745), .B0(N4166), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1419 (.Y(N5109), .A0(N4533), .A1(N4177), .B0(N4363), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1525 (.Y(N4230), .A0(N4896), .A1(N5073), .B0(N5109), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1313 (.Y(N4927), .A0(N4533), .A1(N4599), .B0(N4268), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1252 (.Y(N5032), .A0(N4533), .A1(N4849), .B0(N4592), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1362 (.Y(N4878), .A0(N4896), .A1(N4927), .B0(N5032), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1577 (.Y(N4895), .A0(N4634), .A1(N4230), .B0(N4878), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1064 (.Y(N4172), .A(N4300), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1052 (.Y(N4638), .A0(N13806), .A1(N4300), .B0(N4297), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1096 (.Y(N5119), .A0(N4533), .A1(N4172), .B0(N4638), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I994 (.Y(N4917), .A0(N13795), .A1(N4479), .B0(N13786), .B1(N13766));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1024 (.Y(N4612), .A0(N4533), .A1(N4917), .B0(N4721), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1142 (.Y(N4281), .A0(N4896), .A1(N5119), .B0(N4612), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I838 (.Y(N4855), .A(N4826), .B(N4166));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I898 (.Y(N4933), .A0(N4533), .A1(N5163), .B0(N4855), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I759 (.Y(N4556), .A0(N13791), .A1(N4479), .B0(N4300), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I800 (.Y(N4481), .A0(N4533), .A1(N4556), .B0(N4531), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I946 (.Y(N5110), .A0(N4896), .A1(N4933), .B0(N4481), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1197 (.Y(N4453), .A0(N4634), .A1(N4281), .B0(N5110), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1630 (.Y(N480), .A0(N4911), .A1(N4895), .B0(N4453), .B1(a_man[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1278 (.Y(N4534), .A(N4314), .B(N4297));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1475 (.Y(N4629), .A0(N4533), .A1(N4534), .B0(N5061), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1417 (.Y(N4661), .A0(N4533), .A1(N4918), .B0(N4903), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1523 (.Y(N4807), .A0(N4896), .A1(N4629), .B0(N4661), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1286 (.Y(N4782), .A0(N4314), .A1(N13760), .B0(N4438), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1275 (.Y(N4835), .A0(N4314), .A1(N4166), .B0(N13745), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1311 (.Y(N4480), .A0(N4533), .A1(N4782), .B0(N4835), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1250 (.Y(N4588), .A0(N4948), .A1(N4533), .B0(a_man[19]), .B1(N4431));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1360 (.Y(N4430), .A0(N4896), .A1(N4480), .B0(N4588), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1575 (.Y(N4451), .A0(N4634), .A1(N4807), .B0(N4430), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1051 (.Y(N4986), .A0(N13806), .A1(N13745), .B0(N4438), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1094 (.Y(N4672), .A0(N4533), .A1(N4745), .B0(N4986), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I993 (.Y(N4249), .A(N4280), .B(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5882 (.Y(N4168), .A0(N4533), .A1(N4249), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5889 (.Y(N4850), .A0(N4896), .A1(N4672), .B0(N4168), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I836 (.Y(N4985), .A0(N13806), .A1(N4438), .B0(N4166), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I896 (.Y(N4487), .A0(N4533), .A1(N4435), .B0(N4985), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I757 (.Y(N4915), .A(N13744), .B(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I798 (.Y(N5054), .A0(N4915), .A1(N4533), .B0(a_man[19]), .B1(N4794));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I944 (.Y(N4662), .A0(N4896), .A1(N4487), .B0(N5054), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1195 (.Y(N5027), .A0(N4634), .A1(N4850), .B0(N4662), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1628 (.Y(N478), .A0(N4911), .A1(N4451), .B0(N5027), .B1(a_man[22]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I729 (.Y(N4535), .A(N4314), .B(N4736));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1476 (.Y(N4851), .A0(N4533), .A1(N4535), .B0(N4550), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1418 (.Y(N4883), .A0(N4533), .A1(N4194), .B0(N4918), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1524 (.Y(N5028), .A0(N4896), .A1(N4851), .B0(N4883), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1312 (.Y(N4697), .A0(N4533), .A1(N4411), .B0(N4167), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1251 (.Y(N4810), .A0(N4533), .A1(N4969), .B0(N4939), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1361 (.Y(N4657), .A0(N4896), .A1(N4697), .B0(N4810), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1576 (.Y(N4673), .A0(N4634), .A1(N5028), .B0(N4657), .B1(a_man[21]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I1063 (.Y(N4971), .A(N4438));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1095 (.Y(N4891), .A0(N4533), .A1(N4971), .B0(N13807), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1023 (.Y(N4388), .A0(N4561), .A1(N4533), .B0(a_man[19]), .B1(N4768));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1141 (.Y(N5072), .A0(N4896), .A1(N4891), .B0(N4388), .B1(a_man[20]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I837 (.Y(N4188), .A(N13803), .B(N4869));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I897 (.Y(N4703), .A0(N4533), .A1(N4470), .B0(N4188), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I724 (.Y(N5020), .A0(N4314), .A1(N13745), .B0(N4736), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I799 (.Y(N4259), .A0(N4533), .A1(N5061), .B0(N5020), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I945 (.Y(N4884), .A0(N4896), .A1(N4703), .B0(N4259), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1196 (.Y(N4229), .A0(N4634), .A1(N5072), .B0(N4884), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1629 (.Y(N479), .A0(N4911), .A1(N4673), .B0(N4229), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I16118 (.CO(N8588), .S(N26236), .A(N478), .B(N479));
ADDHX1 inst_cellmath__64_0_I2519 (.CO(N9157), .S(N8994), .A(N480), .B(N8588));
NOR2XL inst_cellmath__63_0_I2192 (.Y(N7475), .A(N3538), .B(N7050));
NOR2XL inst_cellmath__63_0_I2030 (.Y(N7211), .A(N3456), .B(N6952));
NOR2XL inst_cellmath__63_0_I2084 (.Y(N7299), .A(N3611), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2364 (.CO(N6900), .S(N7589), .A(N7475), .B(N7211), .CI(N7299));
NOR2XL inst_cellmath__63_0_I2102 (.Y(N7328), .A(N3702), .B(N7288));
NOR2XL inst_cellmath__63_0_I2156 (.Y(N7414), .A(N3462), .B(N7321));
NOR2XL inst_cellmath__63_0_I2048 (.Y(N7238), .A(N3412), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2363 (.CO(N7394), .S(N7202), .A(N7328), .B(N7414), .CI(N7238));
ADDFX1 inst_cellmath__63_0_I2368 (.CO(N7556), .S(N7365), .A(N7589), .B(N7202), .CI(N7691));
ADDFXL inst_cellmath__63_0_I2371 (.CO(N6946), .S(N7639), .A(N7465), .B(N7365), .CI(N6962));
ADDFX1 inst_cellmath__63_0_I2366 (.CO(N7675), .S(N7481), .A(N6919), .B(N7416), .CI(N7303));
NOR2XL inst_cellmath__63_0_I2012 (.Y(N7183), .A(N3503), .B(N7533));
NOR2XL inst_cellmath__63_0_I1994 (.Y(N7153), .A(N3603), .B(N7304));
NOR2XL inst_cellmath__63_0_I2120 (.Y(N7356), .A(N3399), .B(N7594));
ADDFXL inst_cellmath__63_0_I2362 (.CO(N7011), .S(N7703), .A(N7183), .B(N7153), .CI(N7356));
NAND2X1 inst_cellmath__63_0_I2210 (.Y(N7505), .A(inst_cellmath__48[15]), .B(N7159));
NOR2XL inst_cellmath__63_0_I1958 (.Y(N7100), .A(N7350), .B(N7576));
INVXL inst_cellmath__63_0_I2359 (.Y(N7038), .A(N6885));
ADDFX1 inst_cellmath__63_0_I2360 (.CO(N7621), .S(N7428), .A(N7100), .B(N7505), .CI(N7038));
NOR2XL inst_cellmath__63_0_I2174 (.Y(N7445), .A(N3496), .B(N7627));
NOR2XL inst_cellmath__63_0_I1976 (.Y(N7127), .A(N3142), .B(N6998));
NOR2XL inst_cellmath__63_0_I2138 (.Y(N7384), .A(N3432), .B(N7016));
ADDFX1 inst_cellmath__63_0_I2361 (.CO(N7513), .S(N7317), .A(N7127), .B(N7445), .CI(N7384));
ADDFXL inst_cellmath__63_0_I2367 (.CO(N7171), .S(N6977), .A(N7703), .B(N7428), .CI(N7317));
ADDFX1 inst_cellmath__63_0_I2370 (.CO(N7446), .S(N7250), .A(N7079), .B(N7481), .CI(N6977));
NOR2XL inst_cellmath__63_0_I2066 (.Y(N7266), .A(N3446), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2365 (.CO(N7283), .S(N7095), .A(N7532), .B(N7266), .CI(N7032));
ADDFX1 inst_cellmath__63_0_I2369 (.CO(N7063), .S(N6865), .A(N7095), .B(N7190), .CI(N7575));
ADDFXL inst_cellmath__63_0_I2372 (.CO(N7333), .S(N7142), .A(N6865), .B(N7250), .CI(N7348));
ADDFXL inst_cellmath__63_0_I2373 (.CO(inst_cellmath__63__W0[19]), .S(inst_cellmath__63__W1[18]), .A(N6850), .B(N7639), .CI(N7142));
ADDFXL inst_cellmath__64_0_I2520 (.CO(N8733), .S(N9307), .A(inst_cellmath__63__W0[18]), .B(N8994), .CI(inst_cellmath__63__W1[18]));
ADDFHXL inst_cellmath__64_0_I2525 (.CO(N8866), .S(N8707), .A(inst_cellmath__62__W0[19]), .B(inst_cellmath__62__W1[19]), .CI(N8733));
NOR2XL inst_cellmath__63_0_I2139 (.Y(N6888), .A(N3432), .B(N7594));
NOR2XL inst_cellmath__63_0_I2031 (.Y(N7600), .A(N3456), .B(N7533));
NOR2XL inst_cellmath__63_0_I2103 (.Y(N6835), .A(N3702), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2377 (.CO(N7493), .S(N7298), .A(N6888), .B(N7600), .CI(N6835));
NOR2XL inst_cellmath__63_0_I1977 (.Y(N7515), .A(N3142), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2374 (.CO(N7217), .S(N7028), .A(N6885), .B(N7350), .CI(N7515));
NOR2XL inst_cellmath__63_0_I2175 (.Y(N6945), .A(N3496), .B(N7321));
NOR2XL inst_cellmath__63_0_I2067 (.Y(N7658), .A(N3446), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2378 (.CO(N6992), .S(N7685), .A(N7028), .B(N6945), .CI(N7658));
ADDFX1 inst_cellmath__63_0_I2382 (.CO(N7652), .S(N7459), .A(N7298), .B(N7685), .CI(N7283));
NOR2XL inst_cellmath__63_0_I2085 (.Y(N7686), .A(N3611), .B(N7562));
NOR2XL inst_cellmath__63_0_I2049 (.Y(N7625), .A(N3412), .B(N6952));
ADDFX1 inst_cellmath__63_0_I2379 (.CO(N7376), .S(N7184), .A(N7686), .B(N7625), .CI(N7621));
ADDFXL inst_cellmath__63_0_I2383 (.CO(N7152), .S(N6957), .A(N7675), .B(N7184), .CI(N7171));
ADDFXL inst_cellmath__63_0_I2385 (.CO(N7043), .S(N6847), .A(N7063), .B(N7459), .CI(N6957));
ADDFX1 inst_cellmath__63_0_I2380 (.CO(N6878), .S(N7570), .A(N7011), .B(N7513), .CI(N7394));
NOR2XL inst_cellmath__63_0_I2193 (.Y(N6971), .A(N3538), .B(N7627));
NOR2XL inst_cellmath__63_0_I1995 (.Y(N7540), .A(N3603), .B(N6998));
NAND2XL inst_cellmath__63_0_I2211 (.Y(N7003), .A(inst_cellmath__48[15]), .B(N6855));
ADDFX1 inst_cellmath__63_0_I2375 (.CO(N7606), .S(N7410), .A(N6971), .B(N7540), .CI(N7003));
NOR2X1 inst_cellmath__63_0_I2157 (.Y(N6918), .A(N3462), .B(N7016));
NOR2XL inst_cellmath__63_0_I2013 (.Y(N7568), .A(N3503), .B(N7304));
NOR2XL inst_cellmath__63_0_I2121 (.Y(N6857), .A(N3399), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2376 (.CO(N7108), .S(N6913), .A(N6918), .B(N7568), .CI(N6857));
ADDFX1 inst_cellmath__63_0_I2381 (.CO(N7263), .S(N7074), .A(N6900), .B(N6913), .CI(N7410));
ADDFXL inst_cellmath__63_0_I2384 (.CO(N7538), .S(N7344), .A(N7556), .B(N7570), .CI(N7074));
ADDFXL inst_cellmath__63_0_I2386 (.CO(N7424), .S(N7229), .A(N7344), .B(N7446), .CI(N6946));
ADDFXL inst_cellmath__63_0_I2387 (.CO(inst_cellmath__63__W0[20]), .S(inst_cellmath__63__W1[19]), .A(N7333), .B(N6847), .CI(N7229));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1443 (.Y(N4260), .A0(N4314), .A1(N4869), .B0(N4953), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1387 (.Y(N5131), .A0(N4314), .A1(N4300), .B0(N4280), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1479 (.Y(N4500), .A0(N4533), .A1(N4260), .B0(N5131), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1421 (.Y(N4526), .A0(N4533), .A1(N5096), .B0(N4377), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1527 (.Y(N4676), .A0(N4896), .A1(N4500), .B0(N4526), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1287 (.Y(N5097), .A0(N4314), .A1(N4297), .B0(N4166), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1315 (.Y(N4346), .A0(N5097), .A1(N4533), .B0(a_man[19]), .B1(N4276));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1254 (.Y(N4456), .A0(N4533), .A1(N13788), .B0(N13745), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1364 (.Y(N4306), .A0(N4896), .A1(N4346), .B0(N4456), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1579 (.Y(N4326), .A0(N4634), .A1(N4676), .B0(N4306), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1098 (.Y(N4537), .A0(N4533), .A1(N4162), .B0(N4917), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I980 (.Y(N5040), .A0(N4280), .A1(N13795), .B0(N13760), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1026 (.Y(N5058), .A0(N4533), .A1(N4599), .B0(N5040), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1144 (.Y(N4715), .A0(N4896), .A1(N4537), .B0(N5058), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I900 (.Y(N4353), .A0(N4533), .A1(N4785), .B0(N4435), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I802 (.Y(N4928), .A0(N4533), .A1(N5004), .B0(N4670), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I948 (.Y(N4527), .A0(N4896), .A1(N4353), .B0(N4928), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1199 (.Y(N4898), .A0(N4634), .A1(N4715), .B0(N4527), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1632 (.Y(N482), .A0(N4911), .A1(N4326), .B0(N4898), .B1(a_man[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1478 (.Y(N4282), .A0(N4533), .A1(N5102), .B0(N4307), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1420 (.Y(N4312), .A0(N4533), .A1(N4207), .B0(N4704), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1526 (.Y(N4454), .A0(N4896), .A1(N4282), .B0(N4312), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I987 (.Y(N4818), .A0(N13782), .A1(N4953), .B0(N13745), .B1(N13795));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1314 (.Y(N5146), .A0(N4533), .A1(N5163), .B0(N4818), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1226 (.Y(N4759), .A0(N4314), .A1(N4869), .B0(N4166), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1253 (.Y(N4235), .A0(N4533), .A1(N4759), .B0(N4382), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1363 (.Y(N5104), .A0(N4896), .A1(N5146), .B0(N4235), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1578 (.Y(N5123), .A0(N4634), .A1(N4454), .B0(N5104), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1097 (.Y(N4322), .A0(N4533), .A1(N5020), .B0(N4988), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1025 (.Y(N4836), .A0(N4533), .A1(N4747), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1143 (.Y(N4499), .A0(N4896), .A1(N4322), .B0(N4836), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I867 (.Y(N4558), .A0(N13806), .A1(N13745), .B0(N4280), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I899 (.Y(N5153), .A0(N4533), .A1(N4558), .B0(N4794), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I760 (.Y(N4510), .A0(a_man[17]), .A1(N13795), .B0(N4438), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I801 (.Y(N4698), .A0(N4533), .A1(N4510), .B0(N4981), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I947 (.Y(N4313), .A0(N4896), .A1(N5153), .B0(N4698), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1198 (.Y(N4675), .A0(N4634), .A1(N4499), .B0(N4313), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1631 (.Y(N481), .A0(N4911), .A1(N5123), .B0(N4675), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2523 (.CO(N8970), .S(N8792), .A(N481), .B(N9157));
ADDHX1 inst_cellmath__64_0_I2527 (.CO(N8767), .S(N8605), .A(N482), .B(N8970));
NOR2XL inst_cellmath__63_0_I2176 (.Y(N7331), .A(N3496), .B(N7016));
NOR2XL inst_cellmath__63_0_I2050 (.Y(N7130), .A(N3412), .B(N7533));
NOR2XL inst_cellmath__63_0_I2140 (.Y(N7269), .A(N3432), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2390 (.CO(N7200), .S(N7009), .A(N7331), .B(N7130), .CI(N7269));
NOR2XL inst_cellmath__63_0_I2068 (.Y(N7156), .A(N3446), .B(N6952));
NOR2XL inst_cellmath__63_0_I2158 (.Y(N7302), .A(N3462), .B(N7594));
NOR2XL inst_cellmath__63_0_I2122 (.Y(N7241), .A(N3399), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2391 (.CO(N7587), .S(N7391), .A(N7156), .B(N7302), .CI(N7241));
ADDFX1 inst_cellmath__63_0_I2395 (.CO(N7360), .S(N7166), .A(N7009), .B(N7376), .CI(N7391));
NOR2XL inst_cellmath__63_0_I2086 (.Y(N7185), .A(N3611), .B(N7257));
NOR2XL inst_cellmath__63_0_I2194 (.Y(N7359), .A(N3538), .B(N7321));
NOR2XL inst_cellmath__63_0_I2104 (.Y(N7212), .A(N3702), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2392 (.CO(N7091), .S(N6896), .A(N7185), .B(N7359), .CI(N7212));
NOR2XL inst_cellmath__63_0_I1996 (.Y(N7045), .A(N3603), .B(N7576));
NAND2XL inst_cellmath__63_0_I2212 (.Y(N7386), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[5]));
ADDFX1 inst_cellmath__63_0_I2388 (.CO(N7315), .S(N7123), .A(N7045), .B(N3142), .CI(N7386));
ADDFXL inst_cellmath__63_0_I2393 (.CO(N7477), .S(N7279), .A(N7108), .B(N7606), .CI(N7123));
ADDFXL inst_cellmath__63_0_I2396 (.CO(N6861), .S(N7553), .A(N6878), .B(N6896), .CI(N7279));
ADDFX1 inst_cellmath__63_0_I2398 (.CO(N7634), .S(N7441), .A(N7152), .B(N7166), .CI(N7553));
NOR2XL inst_cellmath__63_0_I2014 (.Y(N7073), .A(N3503), .B(N6998));
NOR2XL inst_cellmath__63_0_I2032 (.Y(N7103), .A(N3456), .B(N7304));
ADDFX1 inst_cellmath__63_0_I2389 (.CO(N7700), .S(N7510), .A(N7217), .B(N7073), .CI(N7103));
ADDFXL inst_cellmath__63_0_I2394 (.CO(N6974), .S(N7669), .A(N7493), .B(N6992), .CI(N7510));
ADDFXL inst_cellmath__63_0_I2397 (.CO(N7247), .S(N7057), .A(N7669), .B(N7263), .CI(N7652));
ADDFXL inst_cellmath__63_0_I2399 (.CO(N7138), .S(N6943), .A(N7057), .B(N7538), .CI(N7043));
ADDFXL inst_cellmath__63_0_I2400 (.CO(inst_cellmath__63__W0[21]), .S(inst_cellmath__63__W1[20]), .A(N7424), .B(N7441), .CI(N6943));
ADDFXL inst_cellmath__64_0_I2528 (.CO(N9098), .S(N8942), .A(N8605), .B(inst_cellmath__63__W0[20]), .CI(inst_cellmath__63__W1[20]));
NOR2XL inst_cellmath__62_0_I1742 (.Y(N6295), .A(N6391), .B(N6286));
NOR2XL inst_cellmath__62_0_I1790 (.Y(N6225), .A(N6347), .B(N6331));
NOR2XL inst_cellmath__62_0_I1766 (.Y(N6428), .A(N6198), .B(N6477));
ADDFX1 inst_cellmath__62_0_I1873 (.CO(N6442), .S(N6365), .A(N6295), .B(N6225), .CI(N6428));
NOR2XL inst_cellmath__62_0_I1754 (.Y(N6360), .A(N6467), .B(N6213));
NOR2XL inst_cellmath__62_0_I1778 (.Y(N6497), .A(N6276), .B(N6404));
ADDFHXL inst_cellmath__62_0_I1874 (.CO(N6253), .S(N6176), .A(N6360), .B(N6497), .CI(N6379));
ADDFHXL inst_cellmath__62_0_I1875 (.CO(N6399), .S(N6323), .A(N6365), .B(N6189), .CI(N6176));
ADDFHXL inst_cellmath__62_0_I1876 (.CO(inst_cellmath__62__W0[21]), .S(inst_cellmath__62__W1[20]), .A(N6486), .B(N6339), .CI(N6323));
ADDFXL inst_cellmath__64_0_I2524 (.CO(N9282), .S(N9128), .A(inst_cellmath__63__W0[19]), .B(N8792), .CI(inst_cellmath__63__W1[19]));
ADDFHXL inst_cellmath__64_0_I2529 (.CO(N8680), .S(N9257), .A(inst_cellmath__62__W0[20]), .B(inst_cellmath__62__W1[20]), .CI(N9282));
ADDFHXL inst_cellmath__64_0_I2530 (.CO(N9007), .S(N8833), .A(N8866), .B(N8942), .CI(N9257));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1480 (.Y(N4716), .A0(N4533), .A1(N4435), .B0(N4308), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1422 (.Y(N4752), .A0(N4533), .A1(N5127), .B0(N4599), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1528 (.Y(N4899), .A0(N4896), .A1(N4716), .B0(N4752), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1280 (.Y(N4404), .A(N4297), .B(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1316 (.Y(N4564), .A0(N4533), .A1(N4404), .B0(N4638), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1227 (.Y(N4409), .A0(N4314), .A1(N4166), .B0(N4479), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1220 (.Y(N5052), .A0(N4314), .A1(N4297), .B0(N13760), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1255 (.Y(N4678), .A0(N4533), .A1(N4409), .B0(N5052), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1365 (.Y(N4522), .A0(N4896), .A1(N4564), .B0(N4678), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1580 (.Y(N4539), .A0(N4634), .A1(N4899), .B0(N4522), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1099 (.Y(N4760), .A0(N4533), .A1(N5064), .B0(N4774), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1027 (.Y(N4264), .A0(N4533), .A1(N4557), .B0(N4786), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1145 (.Y(N4944), .A0(N4896), .A1(N4760), .B0(N4264), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I763 (.Y(N4303), .A0(N13797), .A1(N4869), .B0(N4280), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I901 (.Y(N4574), .A0(N4533), .A1(N4303), .B0(N4948), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I762 (.Y(N4425), .A(N13797), .B(N13745));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I728 (.Y(N4320), .A0(N4314), .A1(N13745), .B0(N4869), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I803 (.Y(N5147), .A0(N4533), .A1(N4425), .B0(N4320), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I949 (.Y(N4753), .A0(N4896), .A1(N4574), .B0(N5147), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1200 (.Y(N5125), .A0(N4634), .A1(N4944), .B0(N4753), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1633 (.Y(N483), .A0(N4911), .A1(N4539), .B0(N5125), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2531 (.CO(N8574), .S(N9172), .A(N483), .B(N8767));
NOR2XL inst_cellmath__63_0_I2051 (.Y(N7518), .A(N3412), .B(N7304));
NAND2XL inst_cellmath__63_0_I2213 (.Y(N6891), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[6]));
NOR2XL inst_cellmath__63_0_I2177 (.Y(N6837), .A(N3496), .B(N7594));
ADDFX1 inst_cellmath__63_0_I2402 (.CO(N7407), .S(N7214), .A(N7518), .B(N6891), .CI(N6837));
NOR2XL inst_cellmath__63_0_I2195 (.Y(N6859), .A(N3538), .B(N7016));
NOR2XL inst_cellmath__63_0_I2069 (.Y(N7542), .A(N3446), .B(N7533));
NOR2XL inst_cellmath__63_0_I2159 (.Y(N7690), .A(N3462), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2403 (.CO(N6910), .S(N7601), .A(N6859), .B(N7542), .CI(N7690));
ADDFX1 inst_cellmath__63_0_I2407 (.CO(N7566), .S(N7372), .A(N7214), .B(N7091), .CI(N7601));
NOR2XL inst_cellmath__63_0_I2141 (.Y(N7661), .A(N3432), .B(N6983));
NOR2XL inst_cellmath__63_0_I2087 (.Y(N7571), .A(N3611), .B(N6952));
NOR2XL inst_cellmath__63_0_I2105 (.Y(N7602), .A(N3702), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2404 (.CO(N7294), .S(N7104), .A(N7661), .B(N7571), .CI(N7602));
ADDFX1 inst_cellmath__63_0_I2408 (.CO(N7071), .S(N6875), .A(N7477), .B(N7104), .CI(N6974));
ADDFX1 inst_cellmath__63_0_I2410 (.CO(N6955), .S(N7648), .A(N6861), .B(N7372), .CI(N6875));
NOR2XL inst_cellmath__63_0_I2123 (.Y(N7630), .A(N3399), .B(N7562));
NOR2XL inst_cellmath__63_0_I2033 (.Y(N7487), .A(N3456), .B(N6998));
NOR2XL inst_cellmath__63_0_I2015 (.Y(N7458), .A(N3503), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2401 (.CO(N7023), .S(N6834), .A(N7487), .B(N7458), .CI(N3603));
ADDFX1 inst_cellmath__63_0_I2405 (.CO(N7682), .S(N7490), .A(N7315), .B(N7630), .CI(N6834));
ADDFX1 inst_cellmath__63_0_I2406 (.CO(N7181), .S(N6987), .A(N7200), .B(N7700), .CI(N7587));
ADDFX1 inst_cellmath__63_0_I2409 (.CO(N7456), .S(N7259), .A(N7360), .B(N7490), .CI(N6987));
ADDFXL inst_cellmath__63_0_I2411 (.CO(N7342), .S(N7150), .A(N7259), .B(N7247), .CI(N7634));
ADDFX1 inst_cellmath__63_0_I2412 (.CO(inst_cellmath__63__W0[22]), .S(inst_cellmath__63__W1[21]), .A(N7138), .B(N7648), .CI(N7150));
ADDFX1 inst_cellmath__64_0_I2532 (.CO(N8913), .S(N8745), .A(inst_cellmath__63__W0[21]), .B(N9172), .CI(inst_cellmath__63__W1[21]));
NOR2XL inst_cellmath__62_0_I1767 (.Y(N6237), .A(N6198), .B(N6213));
NOR2X1 inst_cellmath__62_0_I1779 (.Y(N6305), .A(N6276), .B(N6477));
NOR2X1 inst_cellmath__62_0_I1755 (.Y(N6511), .A(N6467), .B(N6286));
NOR2XL inst_cellmath__62_0_I1791 (.Y(N6371), .A(N6347), .B(N6404));
ADDFXL inst_cellmath__62_0_I1877 (.CO(N6355), .S(N6281), .A(N6305), .B(N6511), .CI(N6371));
ADDFX1 inst_cellmath__62_0_I1878 (.CO(N6502), .S(N6427), .A(N6442), .B(N6237), .CI(N6281));
ADDFX1 inst_cellmath__62_0_I1879 (.CO(inst_cellmath__62__W1[22]), .S(inst_cellmath__62__W1[21]), .A(N6427), .B(N6253), .CI(N6399));
ADDFHXL inst_cellmath__64_0_I2533 (.CO(N9235), .S(N9070), .A(inst_cellmath__62__W1[21]), .B(inst_cellmath__62__W0[21]), .CI(N9098));
ADDFHXL inst_cellmath__64_0_I2534 (.CO(N8805), .S(N8653), .A(N8680), .B(N8745), .CI(N9070));
NAND2X2 inst_cellmath__64_0_I2711 (.Y(N9013), .A(N9007), .B(N8653));
NOR2XL inst_cellmath__62_0_I1688 (.Y(N6498), .A(N6434), .B(N6477));
NOR2XL inst_cellmath__62_0_I1712 (.Y(N6291), .A(N6244), .B(N6331));
NOR2XL inst_cellmath__62_0_I1676 (.Y(N6430), .A(N6359), .B(N6213));
ADDFX1 inst_cellmath__62_0_I1833 (.CO(N6289), .S(N6217), .A(N6498), .B(N6291), .CI(N6430));
ADDFX1 inst_cellmath__62_0_I1843 (.CO(N6413), .S(N6341), .A(N6289), .B(N6423), .CI(N6233));
NOR2XL inst_cellmath__62_0_I1700 (.Y(N6226), .A(N6509), .B(N6404));
NOR2XL inst_cellmath__62_0_I1747 (.Y(N6344), .A(N6467), .B(N6372));
NOR2XL inst_cellmath__62_0_I1735 (.Y(N6278), .A(N6391), .B(N6446));
ADDHX1 inst_cellmath__62_0_I1823 (.CO(N6507), .S(N6432), .A(N6344), .B(N6278));
NAND2BXL inst_noninc_a_cellmath__55_2WWMM_I16171 (.Y(N26407), .AN(N3657), .B(N3739));
XOR2XL inst_noninc_a_cellmath__55_2WWMM_I16180 (.Y(N6492), .A(N3756), .B(N26407));
NOR2XL inst_cellmath__62_0_I1783 (.Y(N6206), .A(N6347), .B(N6492));
NOR2XL inst_cellmath__62_0_I1771 (.Y(N6478), .A(N6276), .B(N6227));
NOR2XL inst_cellmath__62_0_I1723 (.Y(N6211), .A(N6317), .B(N6184));
ADDFX1 inst_cellmath__62_0_I1824 (.CO(N6315), .S(N6242), .A(N6206), .B(N6478), .CI(N6211));
ADDFX1 inst_cellmath__62_0_I1834 (.CO(N6438), .S(N6361), .A(N6226), .B(N6507), .CI(N6315));
NOR2X1 inst_cellmath__62_0_I1711 (.Y(N6484), .A(N6244), .B(N6258));
NOR2XL inst_cellmath__62_0_I1759 (.Y(N6411), .A(N6198), .B(N6298));
NOR2X1 inst_cellmath__62_0_I1699 (.Y(N6416), .A(N6509), .B(N6331));
ADDFX1 inst_cellmath__62_0_I1825 (.CO(N6464), .S(N6389), .A(N6411), .B(N6416), .CI(N6484));
NOR2X1 inst_cellmath__62_0_I1734 (.Y(N6470), .A(N6391), .B(N6372));
NOR2X1 inst_cellmath__62_0_I1722 (.Y(N6403), .A(N6317), .B(N6446));
ADDHXL inst_cellmath__62_0_I1816 (.CO(N6490), .S(N6414), .A(N6403), .B(N6470));
NOR2X1 inst_cellmath__62_0_I1687 (.Y(N6349), .A(N6434), .B(N6404));
NOR2XL inst_cellmath__62_0_I1675 (.Y(N6284), .A(N6359), .B(N6477));
ADDFXL inst_cellmath__62_0_I1826 (.CO(N6273), .S(N6196), .A(N6349), .B(N6490), .CI(N6284));
ADDFXL inst_cellmath__62_0_I1835 (.CO(N6249), .S(N6512), .A(N6464), .B(N6273), .CI(N6262));
ADDFX1 inst_cellmath__62_0_I1844 (.CO(N6223), .S(N6488), .A(N6438), .B(N6380), .CI(N6249));
ADDFHXL inst_cellmath__64_0_I16107 (.CO(N26266), .S(N26253), .A(N6505), .B(N6413), .CI(N6223));
ADDFHXL inst_cellmath__64_0_I16109 (.CO(inst_cellmath__62__W0[18]), .S(N26243), .A(N26266), .B(N6333), .CI(N6480));
NOR2XL inst_cellmath__63_0_I2077 (.Y(N7251), .A(N3611), .B(N7354));
NOR2XL inst_cellmath__63_0_I2095 (.Y(N7277), .A(N3702), .B(N7663));
NOR2XL inst_cellmath__63_0_I1969 (.Y(N7081), .A(N3142), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2271 (.CO(N7281), .S(N7093), .A(N7251), .B(N7277), .CI(N7081));
NOR2XL inst_cellmath__63_0_I1987 (.Y(N7111), .A(N3603), .B(N7594));
NOR2XL inst_cellmath__63_0_I2005 (.Y(N7141), .A(N3503), .B(N7016));
NOR2XL inst_cellmath__63_0_I2059 (.Y(N7222), .A(N3446), .B(N7050));
ADDFX1 inst_cellmath__63_0_I2272 (.CO(N7672), .S(N7479), .A(N7111), .B(N7141), .CI(N7222));
ADDFX1 inst_cellmath__63_0_I2285 (.CO(N7374), .S(N7182), .A(N7281), .B(N7025), .CI(N7672));
ADDFX1 inst_cellmath__63_0_I2299 (.CO(N7474), .S(N7275), .A(N7374), .B(N7508), .CI(N7006));
ADDFXL inst_cellmath__63_0_I2313 (.CO(N7564), .S(N7371), .A(N7102), .B(N7599), .CI(N7474));
ADDFXL inst_cellmath__63_0_I2329 (.CO(N7546), .S(N7353), .A(N7084), .B(N7564), .CI(N7469));
ADDFX1 inst_cellmath__64_0_I16111 (.CO(N26250), .S(N26233), .A(N7546), .B(N7066), .CI(N7452));
ADDFX1 inst_cellmath__64_0_I16119 (.CO(N8928), .S(N26198), .A(N26250), .B(N26236), .CI(N26263));
ADDFXL inst_cellmath__64_0_I2521 (.CO(N9056), .S(N8898), .A(inst_cellmath__62__W0[18]), .B(N8928), .CI(inst_cellmath__62__W1[18]));
ADDFHXL inst_cellmath__64_0_I2526 (.CO(N9197), .S(N9032), .A(N9056), .B(N9128), .CI(N8707));
NAND2X2 inst_cellmath__64_0_I2709 (.Y(N8686), .A(N9197), .B(N8833));
CLKAND2X2 inst_cellmath__64_0_I2780 (.Y(N9092), .A(N9013), .B(N8686));
NOR2XL inst_cellmath__63_0_I2131 (.Y(N7341), .A(N3432), .B(N7310));
NOR2XL inst_cellmath__63_0_I2023 (.Y(N7165), .A(N3456), .B(N7321));
NOR2XL inst_cellmath__63_0_I2113 (.Y(N7312), .A(N3399), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2273 (.CO(N7169), .S(N6975), .A(N7341), .B(N7165), .CI(N7312));
ADDFX1 inst_cellmath__63_0_I2286 (.CO(N6876), .S(N7567), .A(N7408), .B(N7169), .CI(N6911));
NOR2XL inst_cellmath__63_0_I2022 (.Y(N7668), .A(N3456), .B(N7627));
NOR2XL inst_cellmath__63_0_I1932 (.Y(N7524), .A(N6885), .B(N6983));
ADDHX1 inst_cellmath__63_0_I2261 (.CO(N6960), .S(N7654), .A(N7668), .B(N7524));
NOR2XL inst_cellmath__63_0_I1933 (.Y(N7021), .A(N6885), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2274 (.CO(N7554), .S(N7362), .A(N6960), .B(N7021), .CI(N7588));
ADDFX1 inst_cellmath__63_0_I2287 (.CO(N7260), .S(N7072), .A(N7554), .B(N7295), .CI(N7683));
ADDFX1 inst_cellmath__63_0_I2300 (.CO(N6970), .S(N7667), .A(N7389), .B(N6876), .CI(N7260));
ADDFXL inst_cellmath__63_0_I2314 (.CO(N7069), .S(N6873), .A(N6970), .B(N7488), .CI(N6985));
ADDFX1 inst_cellmath__64_0_I16110 (.CO(N26216), .S(N26203), .A(N7069), .B(N6965), .CI(N7353));
INVXL inst_cellmath__64_0_I2511 (.Y(N8840), .A(N478));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1385 (.Y(N4714), .A0(N4314), .A1(a_man[17]), .B0(N13754), .B1(N13788));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1474 (.Y(N4403), .A0(N4533), .A1(N4656), .B0(N4714), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1416 (.Y(N4436), .A0(N4533), .A1(N4250), .B0(N4714), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1522 (.Y(N4583), .A0(N4896), .A1(N4403), .B0(N4436), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1310 (.Y(N4258), .A0(N4533), .A1(N4325), .B0(N4167), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1249 (.Y(N4362), .A0(N4533), .A1(N4745), .B0(N4918), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1359 (.Y(N4210), .A0(N4896), .A1(N4258), .B0(N4362), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1574 (.Y(N4228), .A0(N4634), .A1(N4583), .B0(N4210), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1093 (.Y(N4447), .A0(N4533), .A1(N4290), .B0(N5095), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1021 (.Y(N4965), .A0(N4533), .A1(N4820), .B0(N5159), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1139 (.Y(N4628), .A0(N4896), .A1(N4447), .B0(N4965), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I835 (.Y(N4761), .A0(N13806), .A1(N13745), .B0(N4479), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I895 (.Y(N4265), .A0(N4533), .A1(N4598), .B0(N4761), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I797 (.Y(N4833), .A0(N4533), .A1(N4849), .B0(N4572), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I943 (.Y(N4437), .A0(N4896), .A1(N4265), .B0(N4833), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1194 (.Y(N4806), .A0(N4634), .A1(N4628), .B0(N4437), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1627 (.Y(N477), .A0(N4911), .A1(N4228), .B0(N4806), .B1(a_man[22]));
NOR2XL inst_cellmath__63_0_I1986 (.Y(N7608), .A(N7016), .B(N3603));
NOR2X1 inst_cellmath__63_0_I2040 (.Y(N7694), .A(N3412), .B(N7050));
NOR2XL inst_cellmath__63_0_I1968 (.Y(N7578), .A(N3142), .B(N7594));
ADDFX1 inst_cellmath__63_0_I2263 (.CO(N6848), .S(N7539), .A(N7694), .B(N7608), .CI(N7578));
NOR2XL inst_cellmath__63_0_I2058 (.Y(N6842), .A(N7354), .B(N3446));
NOR2XL inst_cellmath__63_0_I2076 (.Y(N6866), .A(N3611), .B(N7663));
NOR2XL inst_cellmath__63_0_I1950 (.Y(N7548), .A(N7350), .B(N7288));
ADDFXL inst_cellmath__63_0_I2262 (.CO(N7346), .S(N7154), .A(N6842), .B(N6866), .CI(N7548));
NOR2XL inst_cellmath__63_0_I2112 (.Y(N6924), .A(N3399), .B(N7310));
NOR2XL inst_cellmath__63_0_I2004 (.Y(N7637), .A(N3503), .B(N7321));
NOR2XL inst_cellmath__63_0_I2094 (.Y(N6897), .A(N3702), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2264 (.CO(N7232), .S(N7044), .A(N6924), .B(N7637), .CI(N6897));
ADDFX1 inst_cellmath__63_0_I2275 (.CO(N7060), .S(N6863), .A(N6848), .B(N7346), .CI(N7232));
ADDFX1 inst_cellmath__63_0_I2276 (.CO(N7444), .S(N7248), .A(N7479), .B(N7093), .CI(N6975));
ADDFX1 inst_cellmath__63_0_I2288 (.CO(N7650), .S(N7457), .A(N7182), .B(N7060), .CI(N7444));
ADDFX1 inst_cellmath__63_0_I2301 (.CO(N7357), .S(N7164), .A(N7650), .B(N6894), .CI(N7275));
ADDFXL inst_cellmath__63_0_I2315 (.CO(inst_cellmath__63__W0[15]), .S(inst_cellmath__63__W1[14]), .A(N7371), .B(N7357), .CI(N6873));
ADDHX1 inst_cellmath__64_0_I16113 (.CO(N26240), .S(N26222), .A(N477), .B(inst_cellmath__63__W0[15]));
ADDFHXL inst_cellmath__64_0_I16115 (.CO(N26230), .S(N26214), .A(N26216), .B(N8840), .CI(N26240));
NOR2XL inst_cellmath__62_0_I1770 (.Y(N6332), .A(N6276), .B(N6492));
NOR2XL inst_cellmath__62_0_I1758 (.Y(N6266), .A(N6198), .B(N6227));
NOR2XL inst_cellmath__62_0_I1710 (.Y(N6337), .A(N6244), .B(N6184));
ADDFX1 inst_cellmath__62_0_I1817 (.CO(N6296), .S(N6224), .A(N6332), .B(N6266), .CI(N6337));
NOR2XL inst_cellmath__62_0_I1698 (.Y(N6270), .A(N6509), .B(N6258));
NOR2XL inst_cellmath__62_0_I1686 (.Y(N6201), .A(N6434), .B(N6331));
NOR2XL inst_cellmath__62_0_I1746 (.Y(N6195), .A(N6467), .B(N6298));
ADDFX1 inst_cellmath__62_0_I1818 (.CO(N6444), .S(N6370), .A(N6195), .B(N6201), .CI(N6270));
ADDFHXL inst_cellmath__62_0_I1827 (.CO(N6419), .S(N6345), .A(N6432), .B(N6296), .CI(N6444));
ADDFHXL inst_cellmath__62_0_I1836 (.CO(N6396), .S(N6319), .A(N6217), .B(N6408), .CI(N6419));
ADDFXL inst_cellmath__64_0_I16104 (.CO(N26246), .S(N26229), .A(N6190), .B(N6396), .CI(N6341));
ADDFHX1 inst_cellmath__64_0_I16108 (.CO(N26225), .S(N26211), .A(N26246), .B(N26219), .CI(N26253));
ADDFHXL inst_cellmath__64_0_I16120 (.CO(N9246), .S(N26227), .A(N26230), .B(N26225), .CI(N26243));
ADDFHXL inst_cellmath__64_0_I2522 (.CO(N8638), .S(N9223), .A(N9246), .B(N9307), .CI(N8898));
NAND2X2 inst_cellmath__64_0_I2707 (.Y(N9103), .A(N8638), .B(N9032));
NOR2XL inst_cellmath__62_0_I1674 (.Y(N6475), .A(N6359), .B(N6404));
NOR2XL inst_cellmath__62_0_I1721 (.Y(N6257), .A(N6317), .B(N6372));
NOR2XL inst_cellmath__62_0_I1709 (.Y(N6188), .A(N6244), .B(N6446));
ADDHX1 inst_cellmath__62_0_I1810 (.CO(N6279), .S(N6203), .A(N6257), .B(N6188));
ADDFX1 inst_cellmath__62_0_I1819 (.CO(N6256), .S(N6181), .A(N6475), .B(N6279), .CI(N6414));
ADDFX1 inst_cellmath__62_0_I1828 (.CO(N6230), .S(N6496), .A(N6256), .B(N6242), .CI(N6389));
ADDFX1 inst_cellmath__62_0_I1837 (.CO(N6202), .S(N6469), .A(N6230), .B(N6361), .CI(N6512));
ADDFX1 inst_cellmath__64_0_I16105 (.CO(N26206), .S(inst_cellmath__62__W1[15]), .A(N6488), .B(N6202), .CI(N26229));
ADDFXL inst_cellmath__64_0_I16116 (.CO(N26260), .S(N26247), .A(N26214), .B(N26233), .CI(N26206));
ADDFHXL inst_cellmath__64_0_I16121 (.CO(N8820), .S(N8667), .A(N26260), .B(N26198), .CI(N26227));
NAND2X1 inst_cellmath__64_0_I2705 (.Y(N8772), .A(N8820), .B(N9223));
CLKAND2X3 inst_cellmath__64_0_I2778 (.Y(N8859), .A(N9103), .B(N8772));
NAND2X2 inst_cellmath__64_0_I2788 (.Y(N9220), .A(N9092), .B(N8859));
NOR2XL inst_cellmath__62_0_I1685 (.Y(N6393), .A(N6434), .B(N6258));
NOR2XL inst_cellmath__62_0_I1733 (.Y(N6320), .A(N6391), .B(N6298));
NOR2XL inst_cellmath__62_0_I1673 (.Y(N6326), .A(N6359), .B(N6331));
ADDFX1 inst_cellmath__62_0_I1812 (.CO(N6235), .S(N6500), .A(N6393), .B(N6320), .CI(N6326));
NOR2XL inst_cellmath__62_0_I1757 (.Y(N6454), .A(N6198), .B(N6492));
NOR2XL inst_cellmath__62_0_I1745 (.Y(N6387), .A(N6467), .B(N6227));
NOR2XL inst_cellmath__62_0_I1697 (.Y(N6458), .A(N6509), .B(N6184));
ADDFX1 inst_cellmath__62_0_I1811 (.CO(N6425), .S(N6351), .A(N6454), .B(N6387), .CI(N6458));
ADDFX1 inst_cellmath__62_0_I1820 (.CO(N6402), .S(N6328), .A(N6235), .B(N6425), .CI(N6224));
ADDFX1 inst_cellmath__62_0_I1829 (.CO(N6376), .S(N6302), .A(N6402), .B(N6196), .CI(N6345));
ADDFX1 inst_cellmath__64_0_I16103 (.CO(N26213), .S(inst_cellmath__62__W1[14]), .A(N6376), .B(N6319), .CI(N6469));
ADDFX1 inst_cellmath__64_0_I16114 (.CO(N26200), .S(N8720), .A(N26203), .B(N26222), .CI(N26213));
ADDFXL inst_cellmath__64_0_I16117 (.CO(N9019), .S(N8850), .A(N26200), .B(N26211), .CI(N26247));
NAND2X2 inst_cellmath__64_0_I2703 (.Y(N9206), .A(N9019), .B(N8667));
NOR2XL inst_cellmath__63_0_I2003 (.Y(N7249), .A(N3503), .B(N7627));
NOR2XL inst_cellmath__63_0_I2021 (.Y(N7276), .A(N3456), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2253 (.CO(N7413), .S(N7220), .A(N7249), .B(N7276));
NOR2XL inst_cellmath__63_0_I2039 (.Y(N7309), .A(N3412), .B(N7354));
NOR2XL inst_cellmath__63_0_I2057 (.Y(N7338), .A(N3446), .B(N7663));
NOR2XL inst_cellmath__63_0_I1931 (.Y(N7137), .A(N6885), .B(N7288));
ADDFX1 inst_cellmath__63_0_I2254 (.CO(N6916), .S(N7607), .A(N7309), .B(N7338), .CI(N7137));
ADDFX1 inst_cellmath__63_0_I2265 (.CO(N7620), .S(N7427), .A(N7654), .B(N7413), .CI(N6916));
NOR2XL inst_cellmath__63_0_I1949 (.Y(N7161), .A(N7350), .B(N7594));
NOR2XL inst_cellmath__63_0_I1967 (.Y(N7191), .A(N3142), .B(N7016));
NOR2XL inst_cellmath__63_0_I1985 (.Y(N7219), .A(N3603), .B(N7321));
ADDFX1 inst_cellmath__63_0_I2255 (.CO(N7300), .S(N7110), .A(N7161), .B(N7191), .CI(N7219));
ADDFXL inst_cellmath__63_0_I2266 (.CO(N7125), .S(N6927), .A(N7154), .B(N7300), .CI(N7539));
ADDFX1 inst_cellmath__63_0_I2277 (.CO(N6944), .S(N7636), .A(N7362), .B(N7620), .CI(N7125));
ADDFX1 inst_cellmath__63_0_I2289 (.CO(N7151), .S(N6956), .A(N6944), .B(N7567), .CI(N7072));
ADDFX1 inst_cellmath__63_0_I2302 (.CO(inst_cellmath__63__W0[14]), .S(inst_cellmath__63__W1[13]), .A(N7667), .B(N7151), .CI(N7164));
NOR2XL inst_cellmath__62_0_I1708 (.Y(N6378), .A(N6244), .B(N6372));
NOR2XL inst_cellmath__62_0_I1696 (.Y(N6311), .A(N6509), .B(N6446));
ADDHX1 inst_cellmath__62_0_I1805 (.CO(N6218), .S(N6483), .A(N6378), .B(N6311));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I16177 (.Y(N26415), .A(N26407), .B(N3714));
NOR2BX1 inst_noninc_a_cellmath__55_2WWMM_I16178 (.Y(N26417), .AN(N26407), .B(N3756));
NOR3XL inst_noninc_a_cellmath__55_2WWMM_I16179 (.Y(N6241), .A(N6467), .B(N26415), .C(N26417));
NOR2XL inst_cellmath__62_0_I1732 (.Y(N6513), .A(N6391), .B(N6227));
NOR2XL inst_cellmath__62_0_I1684 (.Y(N6246), .A(N6434), .B(N6184));
ADDFX1 inst_cellmath__62_0_I1806 (.CO(N6363), .S(N6290), .A(N6241), .B(N6513), .CI(N6246));
ADDFX1 inst_cellmath__62_0_I1813 (.CO(N6382), .S(N6309), .A(N6203), .B(N6218), .CI(N6363));
ADDFX1 inst_cellmath__62_0_I1821 (.CO(N6210), .S(N6476), .A(N6382), .B(N6370), .CI(N6181));
ADDFX1 inst_cellmath__62_0_I1830 (.CO(inst_cellmath__62__W0[14]), .S(inst_cellmath__62__W1[13]), .A(N6496), .B(N6210), .CI(N6302));
ADDFXL inst_cellmath__64_0_I2506 (.CO(N8657), .S(N9236), .A(inst_cellmath__63__W1[14]), .B(inst_cellmath__63__W0[14]), .CI(inst_cellmath__62__W0[14]));
ADDFXL inst_cellmath__64_0_I16203 (.CO(N9211), .S(N26562), .A(inst_cellmath__62__W1[15]), .B(N8657), .CI(N8720));
NAND2X1 inst_cellmath__64_0_I2701 (.Y(N8873), .A(N9211), .B(N8850));
CLKAND2X2 inst_cellmath__64_0_I2776 (.Y(N8632), .A(N8873), .B(N9206));
NOR2XL inst_cellmath__63_0_I2075 (.Y(N7366), .A(N3611), .B(N7085));
NOR2XL inst_cellmath__63_0_I2093 (.Y(N7392), .A(N3702), .B(N7310));
NOR2XL inst_cellmath__63_0_I1984 (.Y(N6839), .A(N3603), .B(N7627));
NOR2XL inst_cellmath__63_0_I2002 (.Y(N6864), .A(N3503), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2246 (.CO(N7367), .S(N7173), .A(N6839), .B(N6864));
ADDFX1 inst_cellmath__63_0_I2256 (.CO(N7689), .S(N7497), .A(N7366), .B(N7392), .CI(N7367));
NOR2XL inst_cellmath__63_0_I2020 (.Y(N6895), .A(N3456), .B(N7354));
NOR2XL inst_cellmath__63_0_I2038 (.Y(N6922), .A(N3412), .B(N7663));
NOR2XL inst_cellmath__63_0_I1966 (.Y(N7692), .A(N3142), .B(N7321));
ADDFXL inst_cellmath__63_0_I2247 (.CO(N6868), .S(N7559), .A(N6895), .B(N6922), .CI(N7692));
NOR2XL inst_cellmath__63_0_I1930 (.Y(N7632), .A(N6885), .B(N7594));
NOR2XL inst_cellmath__63_0_I1948 (.Y(N7665), .A(N7350), .B(N7016));
NOR2XL inst_cellmath__63_0_I2074 (.Y(N6978), .A(N3611), .B(N7310));
ADDFX1 inst_cellmath__63_0_I2248 (.CO(N7253), .S(N7064), .A(N7632), .B(N7665), .CI(N6978));
ADDFX1 inst_cellmath__63_0_I2257 (.CO(N7187), .S(N6994), .A(N7220), .B(N6868), .CI(N7253));
ADDFX1 inst_cellmath__63_0_I2267 (.CO(N7512), .S(N7316), .A(N7044), .B(N7689), .CI(N7187));
ADDFX1 inst_cellmath__63_0_I2278 (.CO(N7330), .S(N7140), .A(N7512), .B(N6863), .CI(N7248));
ADDFX1 inst_cellmath__63_0_I2290 (.CO(inst_cellmath__63__W0[13]), .S(inst_cellmath__63__W1[12]), .A(N7457), .B(N7330), .CI(N6956));
NOR2XL inst_cellmath__62_0_I1672 (.Y(N6179), .A(N6359), .B(N6258));
NOR2XL inst_cellmath__62_0_I1720 (.Y(N6445), .A(N6317), .B(N6298));
NOR2XL inst_cellmath__62_0_I1695 (.Y(N6503), .A(N6509), .B(N6372));
NOR2X1 inst_cellmath__62_0_I1683 (.Y(N6437), .A(N6434), .B(N6446));
ADDHX1 inst_cellmath__62_0_I1801 (.CO(N6304), .S(N6231), .A(N6437), .B(N6503));
ADDFX1 inst_cellmath__64_0_I16187 (.CO(N6174), .S(N26496), .A(N6179), .B(N6445), .CI(N6304));
ADDFX1 inst_cellmath__62_0_I1814 (.CO(N6192), .S(N6456), .A(N6351), .B(N6174), .CI(N6500));
ADDFX1 inst_cellmath__62_0_I1822 (.CO(inst_cellmath__62__W0[13]), .S(inst_cellmath__62__W1[12]), .A(N6328), .B(N6192), .CI(N6476));
ADDFXL inst_cellmath__64_0_I2504 (.CO(N8747), .S(N8575), .A(inst_cellmath__63__W1[13]), .B(inst_cellmath__63__W0[13]), .CI(inst_cellmath__62__W0[13]));
ADDFXL inst_cellmath__64_0_I16202 (.CO(N26556), .S(N8807), .A(inst_cellmath__62__W1[14]), .B(N8747), .CI(N9236));
AND2XL inst_cellmath__64_0_I16344 (.Y(N26563), .A(N26556), .B(N26562));
NOR2XL inst_cellmath__63_0_I1965 (.Y(N7306), .A(N3142), .B(N7627));
NOR2XL inst_cellmath__63_0_I1983 (.Y(N7335), .A(N3603), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2240 (.CO(N7705), .S(N7514), .A(N7306), .B(N7335));
NOR2XL inst_cellmath__63_0_I2056 (.Y(N6951), .A(N3446), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2249 (.CO(N7641), .S(N7449), .A(N6951), .B(N7705), .CI(N7173));
ADDFX1 inst_cellmath__63_0_I2258 (.CO(N7572), .S(N7378), .A(N7110), .B(N7607), .CI(N7641));
ADDFXL inst_cellmath__63_0_I2268 (.CO(N7010), .S(N7702), .A(N7572), .B(N7427), .CI(N6927));
ADDFX1 inst_cellmath__63_0_I2279 (.CO(inst_cellmath__63__W0[12]), .S(inst_cellmath__63__W1[11]), .A(N7636), .B(N7010), .CI(N7140));
NOR2XL inst_cellmath__62_0_I1731 (.Y(N6362), .A(N6391), .B(N6492));
NOR2XL inst_cellmath__62_0_I1719 (.Y(N6297), .A(N6317), .B(N6227));
NOR2XL inst_cellmath__62_0_I1671 (.Y(N6369), .A(N6359), .B(N6184));
ADDFX1 inst_cellmath__64_0_I16184 (.CO(N26489), .S(N26473), .A(N6362), .B(N6297), .CI(N6369));
ADDFX1 inst_cellmath__64_0_I16188 (.CO(N6321), .S(N26455), .A(N26489), .B(N6483), .CI(N6290));
ADDFX1 inst_cellmath__62_0_I1815 (.CO(inst_cellmath__62__W0[12]), .S(inst_cellmath__62__W1[11]), .A(N6309), .B(N6321), .CI(N6456));
ADDFXL inst_cellmath__64_0_I2502 (.CO(N8835), .S(N8683), .A(inst_cellmath__63__W1[12]), .B(inst_cellmath__63__W0[12]), .CI(inst_cellmath__62__W0[12]));
ADDFXL inst_cellmath__64_0_I2505 (.CO(N9072), .S(N8918), .A(inst_cellmath__62__W1[13]), .B(N8835), .CI(N8575));
NAND2X1 inst_cellmath__64_0_I16204 (.Y(N26548), .A(N9072), .B(N8807));
NOR2XL inst_cellmath__63_0_I2055 (.Y(N7453), .A(N3446), .B(N7310));
NOR2XL inst_cellmath__63_0_I1929 (.Y(N7245), .A(N6885), .B(N7016));
NOR2XL inst_cellmath__63_0_I2037 (.Y(N7420), .A(N3412), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2242 (.CO(N7590), .S(N7396), .A(N7453), .B(N7245), .CI(N7420));
NOR2XL inst_cellmath__63_0_I2001 (.Y(N7363), .A(N3503), .B(N7354));
NOR2XL inst_cellmath__63_0_I2019 (.Y(N7390), .A(N3456), .B(N7663));
NOR2XL inst_cellmath__63_0_I1947 (.Y(N7272), .A(N7350), .B(N7321));
ADDFX1 inst_cellmath__63_0_I2241 (.CO(N7203), .S(N7012), .A(N7363), .B(N7390), .CI(N7272));
ADDFX1 inst_cellmath__63_0_I2250 (.CO(N7145), .S(N6949), .A(N7590), .B(N7203), .CI(N7559));
ADDFXL inst_cellmath__63_0_I2259 (.CO(N7077), .S(N6881), .A(N7145), .B(N7497), .CI(N6994));
ADDFXL inst_cellmath__64_0_I16193 (.CO(inst_cellmath__63__W0[11]), .S(N26468), .A(N7316), .B(N7077), .CI(N7702));
NOR2XL inst_cellmath__62_0_I1718 (.Y(N6491), .A(N6317), .B(N6492));
NOR2XL inst_cellmath__62_0_I1706 (.Y(N6421), .A(N6244), .B(N6227));
NOR2XL inst_cellmath__62_0_I1694 (.Y(N6354), .A(N6509), .B(N6298));
ADDFX1 inst_cellmath__64_0_I16182 (.CO(N26499), .S(N26483), .A(N6491), .B(N6421), .CI(N6354));
NOR2XL inst_cellmath__62_0_I1707 (.Y(N6232), .A(N6244), .B(N6298));
NOR2XL inst_cellmath__62_0_I1682 (.Y(N6288), .A(N6434), .B(N6372));
NOR2XL inst_cellmath__62_0_I1670 (.Y(N6222), .A(N6359), .B(N6446));
ADDHX1 inst_cellmath__62_0_I1798 (.CO(N6197), .S(N6466), .A(N6288), .B(N6222));
ADDFHXL inst_cellmath__64_0_I16185 (.CO(N26449), .S(N26504), .A(N6232), .B(N6197), .CI(N6231));
ADDFX1 inst_cellmath__64_0_I16186 (.CO(N26479), .S(N26464), .A(N26473), .B(N26499), .CI(N26504));
NOR2XL inst_cellmath__63_0_I1946 (.Y(N6892), .A(N7350), .B(N7627));
NOR2XL inst_cellmath__63_0_I1964 (.Y(N6920), .A(N3142), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2235 (.CO(N7543), .S(N7351), .A(N6892), .B(N6920));
NOR2XL inst_cellmath__63_0_I1982 (.Y(N6948), .A(N3603), .B(N7354));
NOR2XL inst_cellmath__63_0_I2000 (.Y(N6976), .A(N3503), .B(N7663));
NOR2XL inst_cellmath__63_0_I1928 (.Y(N6860), .A(N6885), .B(N7321));
ADDFX1 inst_cellmath__63_0_I2236 (.CO(N7047), .S(N6851), .A(N6948), .B(N6976), .CI(N6860));
ADDFX1 inst_cellmath__63_0_I2243 (.CO(N7096), .S(N6901), .A(N7514), .B(N7543), .CI(N7047));
ADDFX1 inst_cellmath__63_0_I2251 (.CO(N7529), .S(N7334), .A(N7096), .B(N7064), .CI(N7449));
ADDFX1 inst_cellmath__64_0_I16192 (.CO(N26452), .S(N26439), .A(N7378), .B(N7529), .CI(N6881));
ADDFXL inst_cellmath__64_0_I16198 (.CO(N9035), .S(N26481), .A(N26452), .B(N26479), .CI(N26468));
ADDFXL inst_cellmath__64_0_I2500 (.CO(N8946), .S(N8770), .A(inst_cellmath__63__W1[11]), .B(inst_cellmath__63__W0[11]), .CI(N9035));
ADDFHXL inst_cellmath__64_0_I2503 (.CO(N9176), .S(N9009), .A(inst_cellmath__62__W1[12]), .B(N8946), .CI(N8683));
AND2XL inst_cellmath__64_0_I2635 (.Y(N8769), .A(N9176), .B(N8918));
ADDFX1 inst_cellmath__64_0_I16189 (.CO(inst_cellmath__62__W0[11]), .S(N26486), .A(N26496), .B(N26449), .CI(N26455));
ADDFXL inst_cellmath__64_0_I2501 (.CO(N9260), .S(N9100), .A(inst_cellmath__62__W1[11]), .B(inst_cellmath__62__W0[11]), .CI(N8770));
NAND2X2 inst_cellmath__64_0_I2633 (.Y(N9199), .A(N9260), .B(N9009));
NOR2XL inst_cellmath__63_0_I1963 (.Y(N7418), .A(N3142), .B(N7354));
NOR2XL inst_cellmath__63_0_I1981 (.Y(N7450), .A(N3603), .B(N7663));
NOR2XL inst_cellmath__63_0_I2017 (.Y(N7509), .A(N3456), .B(N7310));
ADDFX1 inst_cellmath__63_0_I2232 (.CO(N7267), .S(N7080), .A(N7418), .B(N7450), .CI(N7509));
ADDFXL inst_cellmath__63_0_I2238 (.CO(N6931), .S(N7623), .A(N7267), .B(N7351), .CI(N6851));
NOR2XL inst_cellmath__63_0_I2018 (.Y(N7007), .A(N3456), .B(N7085));
NOR2XL inst_cellmath__63_0_I2036 (.Y(N7037), .A(N3412), .B(N7310));
NOR2XL inst_cellmath__63_0_I1927 (.Y(N7358), .A(N6885), .B(N7627));
NOR2XL inst_cellmath__63_0_I1945 (.Y(N7387), .A(N7350), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2231 (.CO(N6886), .S(N7577), .A(N7358), .B(N7387));
ADDFX1 inst_cellmath__63_0_I2237 (.CO(N7430), .S(N7234), .A(N7007), .B(N7037), .CI(N6886));
ADDFX1 inst_cellmath__63_0_I2244 (.CO(N7483), .S(N7284), .A(N7430), .B(N7012), .CI(N7396));
ADDFX1 inst_cellmath__64_0_I16190 (.CO(N26461), .S(inst_cellmath__63__W1[7]), .A(N6931), .B(N6901), .CI(N7284));
NOR2XL inst_cellmath__62_0_I1669 (.Y(N6412), .A(N6359), .B(N6372));
NOR2XL inst_cellmath__62_0_I1705 (.Y(N6275), .A(N6244), .B(N6492));
ADDHX1 inst_cellmath__62_0_I1796 (.CO(N6243), .S(inst_cellmath__62__W0[7]), .A(N6412), .B(N6275));
NOR2XL inst_cellmath__63_0_I1962 (.Y(N7034), .A(N3142), .B(N7663));
NOR2XL inst_cellmath__63_0_I1926 (.Y(N6972), .A(N6885), .B(N7050));
ADDHX1 inst_cellmath__63_0_I2228 (.CO(N7501), .S(N7305), .A(N7034), .B(N6972));
NOR2XL inst_cellmath__63_0_I1999 (.Y(N7480), .A(N3503), .B(N7085));
ADDFXL inst_cellmath__63_0_I2233 (.CO(N7659), .S(N7466), .A(N7501), .B(N7480), .CI(N7577));
ADDFX1 inst_cellmath__63_0_I2239 (.CO(inst_cellmath__63__W0[7]), .S(inst_cellmath__63__W1[6]), .A(N7234), .B(N7659), .CI(N7623));
NOR2XL inst_cellmath__63_0_I1998 (.Y(N7094), .A(N3503), .B(N7310));
NOR2XL inst_cellmath__63_0_I1944 (.Y(N7004), .A(N7350), .B(N7354));
NOR2XL inst_cellmath__63_0_I1980 (.Y(N7065), .A(N3603), .B(N7085));
ADDFX1 inst_cellmath__63_0_I2229 (.CO(N6999), .S(inst_cellmath__63__W0[4]), .A(N7094), .B(N7004), .CI(N7065));
ADDFXL inst_cellmath__63_0_I2234 (.CO(inst_cellmath__63__W0[6]), .S(inst_cellmath__63__W1[5]), .A(N7080), .B(N6999), .CI(N7466));
NOR2XL inst_cellmath__62_0_I1692 (.Y(inst_cellmath__62__W0[6]), .A(N6509), .B(N6492));
NOR2XL inst_cellmath__62_0_I1679 (.Y(inst_cellmath__62__W1[5]), .A(N6434), .B(N6492));
NOR2XL inst_cellmath__62_0_I1667 (.Y(inst_cellmath__62__W0[5]), .A(N6359), .B(N6227));
ADDHX1 inst_cellmath__64_0_I2488 (.CO(N8760), .S(N8593), .A(inst_cellmath__62__W1[5]), .B(inst_cellmath__62__W0[5]));
ADDFX1 inst_cellmath__64_0_I2490 (.CO(N8671), .S(N9252), .A(inst_cellmath__63__W0[6]), .B(inst_cellmath__62__W0[6]), .CI(N8760));
ADDFX1 inst_cellmath__64_0_I16194 (.CO(N26444), .S(N9162), .A(inst_cellmath__62__W0[7]), .B(inst_cellmath__63__W0[7]), .CI(N8671));
ADDFX1 inst_cellmath__64_0_I16195 (.CO(N26474), .S(N9061), .A(N26483), .B(N26461), .CI(N26444));
NOR2XL inst_cellmath__62_0_I1681 (.Y(N6479), .A(N6434), .B(N6298));
NOR2XL inst_cellmath__62_0_I1693 (.Y(N6207), .A(N6509), .B(N6227));
NOR2XL inst_cellmath__62_0_I1680 (.Y(N6334), .A(N6434), .B(N6227));
NOR2XL inst_cellmath__62_0_I1668 (.Y(N6268), .A(N6359), .B(N6298));
ADDHX1 inst_cellmath__62_0_I1795 (.CO(N6433), .S(inst_cellmath__62__W1[6]), .A(N6334), .B(N6268));
ADDFX1 inst_cellmath__62_0_I1797 (.CO(N6390), .S(inst_cellmath__62__W1[7]), .A(N6479), .B(N6207), .CI(N6433));
ADDFX1 inst_cellmath__64_0_I16183 (.CO(N26458), .S(inst_cellmath__62__W1[8]), .A(N6243), .B(N6466), .CI(N6390));
ADDFX1 inst_cellmath__64_0_I16191 (.CO(N26493), .S(inst_cellmath__63__W1[8]), .A(N6949), .B(N7483), .CI(N7334));
ADDFXL inst_cellmath__64_0_I16196 (.CO(N26436), .S(N26490), .A(N26458), .B(N26493), .CI(N26439));
ADDFXL inst_cellmath__64_0_I16197 (.CO(N8711), .S(N9285), .A(N26464), .B(N26474), .CI(N26490));
ADDFX1 inst_cellmath__64_0_I16199 (.CO(N8607), .S(N9203), .A(N26436), .B(N26481), .CI(N26486));
NAND2X1 inst_cellmath__64_0_I16200 (.Y(N9283), .A(N8711), .B(N9203));
NOR2XL inst_cellmath__62_0_I1666 (.Y(inst_cellmath__62__W0[4]), .A(N6359), .B(N6492));
ADDHX1 inst_cellmath__64_0_I2487 (.CO(N9190), .S(N9024), .A(inst_cellmath__62__W0[4]), .B(inst_cellmath__63__W0[4]));
NOR2XL inst_cellmath__63_0_I1943 (.Y(N7506), .A(N7350), .B(N7663));
NOR2XL inst_cellmath__63_0_I1925 (.Y(N7476), .A(N6885), .B(N7354));
ADDHX1 inst_cellmath__63_0_I2226 (.CO(N7612), .S(N7417), .A(N7506), .B(N7476));
NOR2XL inst_cellmath__63_0_I1961 (.Y(N7534), .A(N3142), .B(N7085));
NOR2XL inst_cellmath__63_0_I1979 (.Y(N7558), .A(N3603), .B(N7310));
ADDFX1 inst_cellmath__63_0_I2227 (.CO(N7115), .S(inst_cellmath__63__W1[3]), .A(N7534), .B(N7558), .CI(N7417));
ADDFX1 inst_cellmath__63_0_I2230 (.CO(inst_cellmath__63__W0[5]), .S(inst_cellmath__63__W1[4]), .A(N7305), .B(N7612), .CI(N7115));
ADDFX1 inst_cellmath__64_0_I2489 (.CO(N9088), .S(N8934), .A(N9190), .B(inst_cellmath__63__W0[5]), .CI(inst_cellmath__63__W1[5]));
ADDFX1 inst_cellmath__64_0_I2491 (.CO(N8999), .S(N8824), .A(inst_cellmath__62__W1[6]), .B(inst_cellmath__63__W1[6]), .CI(N9088));
ADDFXL inst_cellmath__64_0_I2493 (.CO(N8901), .S(N8738), .A(inst_cellmath__62__W1[7]), .B(inst_cellmath__63__W1[7]), .CI(N8999));
ADDFXL inst_cellmath__64_0_I2495 (.CO(N8797), .S(N8642), .A(inst_cellmath__62__W1[8]), .B(inst_cellmath__63__W1[8]), .CI(N8901));
AND2X1 inst_cellmath__64_0_I2627 (.Y(N8971), .A(N9285), .B(N8797));
AND2XL inst_cellmath__64_0_I2623 (.Y(N9059), .A(N9162), .B(N8738));
NAND2XL inst_cellmath__64_0_I2621 (.Y(N8734), .A(N9252), .B(N8824));
AND2XL inst_cellmath__64_0_I2619 (.Y(N9158), .A(N8593), .B(N8934));
NAND2XL inst_cellmath__64_0_I2617 (.Y(N8822), .A(inst_cellmath__63__W1[4]), .B(N9024));
NOR2XL inst_cellmath__63_0_I1924 (.Y(N7089), .A(N6885), .B(N7663));
NOR2XL inst_cellmath__63_0_I1960 (.Y(N7148), .A(N3142), .B(N7310));
ADDHX1 inst_cellmath__63_0_I2225 (.CO(inst_cellmath__63__W0[3]), .S(inst_cellmath__63__W1[2]), .A(N7089), .B(N7148));
AND2XL inst_cellmath__64_0_I2615 (.Y(N9248), .A(inst_cellmath__63__W1[3]), .B(inst_cellmath__63__W0[3]));
NOR2XL inst_cellmath__63_0_I1942 (.Y(inst_cellmath__63__W0[2]), .A(N7350), .B(N7085));
NAND2XL inst_cellmath__64_0_I2613 (.Y(N8931), .A(inst_cellmath__63__W1[2]), .B(inst_cellmath__63__W0[2]));
OR4X1 inst_cellmath__64_0_I16301 (.Y(N8655), .A(N7350), .B(N6885), .C(N7310), .D(N7085));
NOR2XL inst_cellmath__64_0_I2612 (.Y(N8756), .A(inst_cellmath__63__W1[2]), .B(inst_cellmath__63__W0[2]));
AOI21XL inst_cellmath__64_0_I2642 (.Y(N9210), .A0(N8931), .A1(N8655), .B0(N8756));
OAI22XL inst_cellmath__64_0_I5924 (.Y(N8926), .A0(N9248), .A1(N9210), .B0(inst_cellmath__63__W1[3]), .B1(inst_cellmath__63__W0[3]));
NOR2XL inst_cellmath__64_0_I2616 (.Y(N8668), .A(inst_cellmath__63__W1[4]), .B(N9024));
AOI21XL inst_cellmath__64_0_I2646 (.Y(N8636), .A0(N8822), .A1(N8926), .B0(N8668));
OAI22XL inst_cellmath__64_0_I5925 (.Y(N9006), .A0(N9158), .A1(N8636), .B0(N8593), .B1(N8934));
NOR2XL inst_cellmath__64_0_I2620 (.Y(N8562), .A(N9252), .B(N8824));
AOI21XL inst_cellmath__64_0_I2650 (.Y(N8617), .A0(N8734), .A1(N9006), .B0(N8562));
OAI22XL inst_cellmath__64_0_I5926 (.Y(N8892), .A0(N9059), .A1(N8617), .B0(N9162), .B1(N8738));
NAND2XL inst_cellmath__64_0_I2625 (.Y(N8639), .A(N9061), .B(N8642));
AOI2BB2X1 inst_cellmath__64_0_I5927 (.Y(N9165), .A0N(N9061), .A1N(N8642), .B0(N8892), .B1(N8639));
OR2XL inst_cellmath__64_0_I2626 (.Y(N8795), .A(N8797), .B(N9285));
OAI21X1 inst_cellmath__64_0_I2657 (.Y(N8579), .A0(N8971), .A1(N9165), .B0(N8795));
NOR2XL inst_cellmath__64_0_I2628 (.Y(N9130), .A(N8711), .B(N9203));
AOI21X1 inst_cellmath__64_0_I2658 (.Y(N8762), .A0(N9283), .A1(N8579), .B0(N9130));
AND2XL inst_cellmath__64_0_I2631 (.Y(N8868), .A(N8607), .B(N9100));
OR2XL inst_cellmath__64_0_I2630 (.Y(N8708), .A(N8607), .B(N9100));
OAI21X2 inst_cellmath__64_0_I2661 (.Y(N8836), .A0(N8762), .A1(N8868), .B0(N8708));
NOR2X1 inst_cellmath__64_0_I2632 (.Y(N9034), .A(N9260), .B(N9009));
AOI21X2 inst_cellmath__64_0_I2662 (.Y(N8930), .A0(N9199), .A1(N8836), .B0(N9034));
OR2XL inst_cellmath__64_0_I2634 (.Y(N8606), .A(N9176), .B(N8918));
OAI21X2 inst_cellmath__64_0_I16205 (.Y(N26553), .A0(N8769), .A1(N8930), .B0(N8606));
NOR2XL inst_cellmath__64_0_I2636 (.Y(N8944), .A(N9072), .B(N8807));
AOI21X2 inst_cellmath__64_0_I16211 (.Y(N26561), .A0(N26548), .A1(N26553), .B0(N8944));
OR2XL inst_cellmath__64_0_I16312 (.Y(N26565), .A(N26556), .B(N26562));
OAI21X4 inst_cellmath__64_0_I16212 (.Y(N8727), .A0(N26563), .A1(N26561), .B0(N26565));
NOR2X2 inst_cellmath__64_0_I2700 (.Y(N8715), .A(N9211), .B(N8850));
NOR2X1 inst_cellmath__64_0_I16122 (.Y(N9038), .A(N9019), .B(N8667));
AOI21X2 inst_cellmath__64_0_I2747 (.Y(N9288), .A0(N8715), .A1(N9206), .B0(N9038));
INVX3 inst_cellmath__64_0_I2775 (.Y(N9217), .A(N9288));
AOI21X4 inst_cellmath__64_0_I2784 (.Y(N9154), .A0(N8727), .A1(N8632), .B0(N9217));
NOR2X1 inst_cellmath__64_0_I2704 (.Y(N8610), .A(N8820), .B(N9223));
NOR2XL inst_cellmath__64_0_I2706 (.Y(N8949), .A(N8638), .B(N9032));
AOI21X2 inst_cellmath__64_0_I2748 (.Y(N9202), .A0(N8610), .A1(N9103), .B0(N8949));
INVX3 inst_cellmath__64_0_I2777 (.Y(N9122), .A(N9202));
NOR2X2 inst_cellmath__64_0_I2708 (.Y(N9262), .A(N9197), .B(N8833));
NOR2XL inst_cellmath__64_0_I2710 (.Y(N8839), .A(N9007), .B(N8653));
AOI21X2 inst_cellmath__64_0_I5774 (.Y(N13738), .A0(N9013), .A1(N9262), .B0(N8839));
INVX2 inst_cellmath__64_0_I5775 (.Y(N8598), .A(N13738));
AOI21X4 inst_cellmath__64_0_I2787 (.Y(N9053), .A0(N9092), .A1(N9122), .B0(N8598));
OAI21X4 cynw_cm_float_rcp_I16259 (.Y(N8674), .A0(N9220), .A1(N9154), .B0(N9053));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1493 (.Y(N4994), .A0(N4533), .A1(N13752), .B0(N4875), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1435 (.Y(N4585), .A0(N4533), .A1(N4154), .B0(N4457), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1541 (.Y(N4728), .A0(N4896), .A1(N4994), .B0(N4585), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1329 (.Y(N4400), .A0(N4533), .A1(N5108), .B0(N4879), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1267 (.Y(N4158), .A0(a_man[17]), .A1(N4533), .B0(N4151), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1378 (.Y(N4358), .A0(N4896), .A1(N4400), .B0(N4158), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1593 (.Y(N4369), .A0(N4634), .A1(N4728), .B0(N4358), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1112 (.Y(N4594), .A0(N4533), .A1(N5046), .B0(N4958), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1040 (.Y(N5117), .A0(N4276), .A1(N4533), .B0(a_man[19]), .B1(N5061));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1158 (.Y(N4770), .A0(N4896), .A1(N4594), .B0(N5117), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I914 (.Y(N4631), .A0(N4290), .A1(N4533), .B0(a_man[19]), .B1(N4276));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I816 (.Y(N4627), .A0(N4533), .A1(N4252), .B0(N13797), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I962 (.Y(N4586), .A0(N4896), .A1(N4631), .B0(N4627), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1213 (.Y(N4954), .A0(N4634), .A1(N4770), .B0(N4586), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1646 (.Y(N496), .A0(N4911), .A1(N4369), .B0(N4954), .B1(a_man[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1492 (.Y(N4334), .A(N4533), .B(N4290));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1434 (.Y(N4360), .A0(N4533), .A1(N4739), .B0(N5108), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1540 (.Y(N4508), .A0(N4896), .A1(N4334), .B0(N4360), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1328 (.Y(N4180), .A0(N4533), .A1(N5127), .B0(N4307), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1266 (.Y(N4957), .A0(N4533), .A1(N13754), .B0(N4818), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1377 (.Y(N5157), .A0(N4896), .A1(N4180), .B0(N4957), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1592 (.Y(N4152), .A0(N4634), .A1(N4508), .B0(N5157), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1111 (.Y(N4367), .A0(N4533), .A1(N4969), .B0(N5140), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1039 (.Y(N4890), .A0(N4533), .A1(N4207), .B0(N4177), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1157 (.Y(N4546), .A0(N4896), .A1(N4367), .B0(N4890), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I873 (.Y(N4935), .A0(a_man[17]), .A1(N13803), .B0(N4953), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I851 (.Y(N4777), .A0(N13760), .A1(N13803), .B0(N13764), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I913 (.Y(N4405), .A0(N4533), .A1(N4935), .B0(N4777), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I815 (.Y(N4401), .A0(N4533), .A1(N5022), .B0(N13760), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I961 (.Y(N4361), .A0(N4896), .A1(N4405), .B0(N4401), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1212 (.Y(N4727), .A0(N4634), .A1(N4546), .B0(N4361), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1645 (.Y(N495), .A0(N4911), .A1(N4152), .B0(N4727), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2581 (.CO(N9192), .S(N9026), .A(inst_cellmath__48[15]), .B(N495));
OR2XL hap1_A_I6066 (.Y(N8567), .A(N496), .B(N9192));
NAND2XL inst_cellmath__64_0_I2739 (.Y(N9090), .A(N8976), .B(N8567));
XNOR2X1 hap1_A_I6065 (.Y(N9164), .A(N496), .B(N9192));
NAND2XL inst_cellmath__63_0_I2223 (.Y(N7205), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[16]));
NOR2XL inst_cellmath__63_0_I2205 (.Y(N7179), .A(N3538), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2476 (.CO(N7656), .S(N7463), .A(N7205), .B(N7179), .CI(N3496));
NAND2XL inst_cellmath__63_0_I2224 (.Y(N7595), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[17]));
ADDFX1 inst_cellmath__63_0_I2478 (.CO(inst_cellmath__63__W1[33]), .S(inst_cellmath__63__W0[32]), .A(N7656), .B(N7595), .CI(N3538));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1491 (.Y(N5133), .A0(N4533), .A1(N5088), .B0(N4777), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1433 (.Y(N5160), .A0(N4533), .A1(N13754), .B0(N4457), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1539 (.Y(N4292), .A0(N4896), .A1(N5133), .B0(N5160), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1327 (.Y(N4980), .A0(N4533), .A1(N4576), .B0(N13788), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1376 (.Y(N4938), .A0(N4896), .A1(N4980), .B0(N4505), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1591 (.Y(N4952), .A0(N4634), .A1(N4292), .B0(N4938), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1110 (.Y(N4149), .A0(N4533), .A1(N4706), .B0(N5101), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1038 (.Y(N4669), .A0(N5062), .A1(N4533), .B0(N4656), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1156 (.Y(N4333), .A0(N4896), .A1(N4149), .B0(N4669), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I912 (.Y(N4183), .A0(N4431), .A1(N4533), .B0(a_man[19]), .B1(N4805));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I814 (.Y(N4181), .A0(N4533), .A1(N4377), .B0(N13744), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I960 (.Y(N5161), .A0(N4896), .A1(N4183), .B0(N4181), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1211 (.Y(N4507), .A0(N4634), .A1(N4333), .B0(N5161), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1644 (.Y(N494), .A0(N4911), .A1(N4952), .B0(N4507), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2577 (.CO(N8631), .S(N9218), .A(N494), .B(inst_cellmath__63__W0[32]));
ADDFX1 inst_cellmath__64_0_I2582 (.CO(N8764), .S(N8597), .A(N9026), .B(inst_cellmath__63__W1[33]), .CI(N8631));
NAND2XL inst_cellmath__64_0_I2737 (.Y(N8759), .A(N9164), .B(N8764));
NAND2XL inst_cellmath__64_0_I2768 (.Y(N8969), .A(N9090), .B(N8759));
NOR2XL inst_cellmath__63_0_I2186 (.Y(N7651), .A(N3496), .B(N7576));
NAND2XL inst_cellmath__63_0_I2222 (.Y(N7710), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[15]));
ADDFX1 inst_cellmath__63_0_I2473 (.CO(N7380), .S(N7188), .A(N7651), .B(N3462), .CI(N7710));
NOR2XL inst_cellmath__63_0_I2167 (.Y(N7233), .A(N3462), .B(N7576));
NAND2XL inst_cellmath__63_0_I2221 (.Y(N7322), .A(inst_cellmath__48[15]), .B(N7339));
ADDFX1 inst_cellmath__63_0_I2469 (.CO(N7609), .S(N7415), .A(N7322), .B(N7233), .CI(N3432));
NOR2XL inst_cellmath__63_0_I2204 (.Y(N7680), .A(N3538), .B(N6998));
ADDFX1 inst_cellmath__63_0_I2474 (.CO(N6882), .S(N7573), .A(N7609), .B(N7680), .CI(N7188));
ADDFX1 inst_cellmath__63_0_I2477 (.CO(inst_cellmath__63__W1[32]), .S(inst_cellmath__63__W0[31]), .A(N7463), .B(N7380), .CI(N6882));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1445 (.Y(N5148), .A0(N4314), .A1(N13754), .B0(N13760), .B1(N13772));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1490 (.Y(N4906), .A0(N4533), .A1(N4534), .B0(N5148), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1432 (.Y(N4941), .A0(N4533), .A1(N4759), .B0(N4935), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1538 (.Y(N5083), .A0(N4896), .A1(N4906), .B0(N4941), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1326 (.Y(N4754), .A0(N4533), .A1(N4969), .B0(N4786), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1265 (.Y(N4862), .A(N4706), .B(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1375 (.Y(N4709), .A0(N4896), .A1(N4754), .B0(N4862), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1590 (.Y(N4724), .A0(N4634), .A1(N5083), .B0(N4709), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1109 (.Y(N4947), .A0(N4656), .A1(N4533), .B0(a_man[19]), .B1(N4431));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1037 (.Y(N4445), .A0(N4533), .A1(N4969), .B0(N4177), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1155 (.Y(N5132), .A0(N4896), .A1(N4947), .B0(N4445), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I911 (.Y(N4982), .A0(N4533), .A1(N13760), .B0(N5061), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I959 (.Y(N4942), .A0(N4896), .A1(N4982), .B0(N4529), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1210 (.Y(N4291), .A0(N4634), .A1(N5132), .B0(N4942), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1643 (.Y(N493), .A0(N4911), .A1(N4724), .B0(N4291), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2573 (.CO(N8814), .S(N8662), .A(N493), .B(inst_cellmath__63__W0[31]));
ADDFX1 inst_cellmath__64_0_I16081 (.CO(N8963), .S(N26158), .A(inst_cellmath__63__W1[32]), .B(N9218), .CI(N8814));
NAND2XL inst_cellmath__64_0_I2735 (.Y(N9189), .A(N8597), .B(N8963));
NOR2XL inst_cellmath__63_0_I2203 (.Y(N7293), .A(N3538), .B(N7304));
NOR2XL inst_cellmath__63_0_I2185 (.Y(N7261), .A(N3496), .B(N6998));
NOR2XL inst_cellmath__63_0_I2166 (.Y(N6849), .A(N3462), .B(N6998));
NOR2XL inst_cellmath__63_0_I2148 (.Y(N7707), .A(N3432), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2464 (.CO(N7451), .S(N7254), .A(N6849), .B(N7707), .CI(N3399));
ADDFX1 inst_cellmath__63_0_I2470 (.CO(N7112), .S(N6917), .A(N7293), .B(N7261), .CI(N7451));
NOR2XL inst_cellmath__63_0_I2184 (.Y(N6877), .A(N3496), .B(N7304));
NAND2XL inst_cellmath__63_0_I2220 (.Y(N6935), .A(inst_cellmath__48[15]), .B(N7645));
NOR2XL inst_cellmath__63_0_I2202 (.Y(N6908), .A(N3538), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2465 (.CO(N6950), .S(N7642), .A(N6877), .B(N6935), .CI(N6908));
ADDFX1 inst_cellmath__63_0_I2471 (.CO(N7498), .S(N7301), .A(N6950), .B(N7415), .CI(N6917));
ADDFX1 inst_cellmath__63_0_I2475 (.CO(inst_cellmath__63__W1[31]), .S(inst_cellmath__63__W0[30]), .A(N7573), .B(N7112), .CI(N7498));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1449 (.Y(N4285), .A0(N4314), .A1(N4166), .B0(N13766), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1489 (.Y(N4681), .A0(N4533), .A1(N4285), .B0(N4835), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1431 (.Y(N4711), .A0(N4533), .A1(N5064), .B0(N5087), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1537 (.Y(N4860), .A0(N4896), .A1(N4681), .B0(N4711), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1325 (.Y(N4528), .A0(N4533), .A1(N4404), .B0(N4818), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1264 (.Y(N4643), .A0(N4533), .A1(N4968), .B0(N5022), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1374 (.Y(N4492), .A0(N4896), .A1(N4528), .B0(N4643), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1589 (.Y(N4506), .A0(N4634), .A1(N4860), .B0(N4492), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1054 (.Y(N4245), .A(N13806), .B(N4869));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1108 (.Y(N4722), .A0(N4533), .A1(N4207), .B0(N4245), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1036 (.Y(N4223), .A0(N4533), .A1(N5141), .B0(N5022), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1154 (.Y(N4905), .A0(N4896), .A1(N4722), .B0(N4223), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I910 (.Y(N4756), .A0(N4533), .A1(N13752), .B0(N4177), .B1(a_man[19]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I812 (.Y(N5112), .A(N4533), .B(N4615));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I958 (.Y(N4712), .A0(N4896), .A1(N4756), .B0(N5112), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1209 (.Y(N5082), .A0(N4634), .A1(N4905), .B0(N4712), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1642 (.Y(N492), .A0(N4911), .A1(N4506), .B0(N5082), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2569 (.CO(N9014), .S(N8843), .A(N492), .B(inst_cellmath__63__W0[30]));
ADDFX1 inst_cellmath__64_0_I16080 (.CO(N26147), .S(N8988), .A(inst_cellmath__63__W1[31]), .B(N8662), .CI(N9014));
NAND2XL inst_cellmath__64_0_I16083 (.Y(N8857), .A(N26158), .B(N26147));
NAND2XL inst_cellmath__64_0_I2765 (.Y(N9057), .A(N9189), .B(N8857));
NOR2XL inst_cellmath__64_0_I2770 (.Y(N8768), .A(N8969), .B(N9057));
NOR2XL inst_cellmath__63_0_I2147 (.Y(N7319), .A(N3432), .B(N6998));
NOR2XL inst_cellmath__63_0_I2129 (.Y(N7290), .A(N3399), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2458 (.CO(N6902), .S(N7591), .A(N7319), .B(N7290), .CI(N3702));
NOR2XL inst_cellmath__63_0_I2165 (.Y(N7347), .A(N3462), .B(N7304));
NAND2XL inst_cellmath__63_0_I2219 (.Y(N7435), .A(inst_cellmath__48[15]), .B(N7067));
NOR2XL inst_cellmath__63_0_I2183 (.Y(N7375), .A(N3496), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2459 (.CO(N7285), .S(N7097), .A(N7347), .B(N7435), .CI(N7375));
ADDFX1 inst_cellmath__63_0_I2466 (.CO(N7336), .S(N7147), .A(N7254), .B(N6902), .CI(N7285));
NOR2XL inst_cellmath__63_0_I2128 (.Y(N6905), .A(N3399), .B(N6998));
NOR2XL inst_cellmath__63_0_I2110 (.Y(N6874), .A(N3702), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2451 (.CO(N6853), .S(N7544), .A(N6905), .B(N6874), .CI(N3611));
NOR2XL inst_cellmath__63_0_I2201 (.Y(N7405), .A(N3538), .B(N6952));
ADDFX1 inst_cellmath__63_0_I2460 (.CO(N7676), .S(N7484), .A(N6853), .B(N7405), .CI(N7591));
ADDFX1 inst_cellmath__63_0_I2467 (.CO(N6840), .S(N7530), .A(N7676), .B(N7642), .CI(N7147));
ADDFX1 inst_cellmath__63_0_I2472 (.CO(inst_cellmath__63__W1[30]), .S(inst_cellmath__63__W0[29]), .A(N7301), .B(N7336), .CI(N6840));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1444 (.Y(N4482), .A(N4314), .B(N13766));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1488 (.Y(N4461), .A0(N4533), .A1(N4308), .B0(N4482), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1430 (.Y(N4497), .A0(N4533), .A1(N5131), .B0(N4652), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1536 (.Y(N4641), .A0(N4896), .A1(N4461), .B0(N4497), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1324 (.Y(N4315), .A0(N4533), .A1(N4519), .B0(N4404), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1263 (.Y(N4416), .A0(N4533), .A1(N4894), .B0(N4818), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1373 (.Y(N4272), .A0(N4896), .A1(N4315), .B0(N4416), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1588 (.Y(N4288), .A0(N4634), .A1(N4641), .B0(N4272), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1107 (.Y(N4504), .A0(N4533), .A1(N4249), .B0(N4747), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1035 (.Y(N5019), .A0(N4533), .A1(N4519), .B0(N4818), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1153 (.Y(N4680), .A0(N4896), .A1(N4504), .B0(N5019), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I909 (.Y(N4536), .A0(N4849), .A1(N4533), .B0(N4939), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I811 (.Y(N4886), .A0(N4533), .A1(N4390), .B0(N4849), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I957 (.Y(N4498), .A0(N4896), .A1(N4536), .B0(N4886), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1208 (.Y(N4859), .A0(N4634), .A1(N4680), .B0(N4498), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1641 (.Y(N491), .A0(N4911), .A1(N4288), .B0(N4859), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2565 (.CO(N9207), .S(N9039), .A(N491), .B(inst_cellmath__63__W0[29]));
ADDFX1 inst_cellmath__64_0_I2570 (.CO(N8581), .S(N9180), .A(N8843), .B(inst_cellmath__63__W1[30]), .CI(N9207));
NAND2XL inst_cellmath__64_0_I2731 (.Y(N9273), .A(N8988), .B(N8581));
NOR2XL inst_cellmath__63_0_I2127 (.Y(N7402), .A(N3399), .B(N7304));
NAND2XL inst_cellmath__63_0_I2217 (.Y(N7547), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[10]));
NOR2XL inst_cellmath__63_0_I2145 (.Y(N7432), .A(N3432), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2444 (.CO(N7693), .S(N7502), .A(N7402), .B(N7547), .CI(N7432));
NOR2XL inst_cellmath__63_0_I2181 (.Y(N7492), .A(N3496), .B(N7257));
NOR2XL inst_cellmath__63_0_I2163 (.Y(N7464), .A(N3462), .B(N6952));
NOR2XL inst_cellmath__63_0_I2199 (.Y(N7523), .A(N3538), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2445 (.CO(N7192), .S(N7000), .A(N7492), .B(N7464), .CI(N7523));
ADDFX1 inst_cellmath__63_0_I2454 (.CO(N7128), .S(N6932), .A(N7693), .B(N7544), .CI(N7192));
NOR2XL inst_cellmath__63_0_I2200 (.Y(N7022), .A(N3538), .B(N7257));
NOR2XL inst_cellmath__63_0_I2182 (.Y(N6990), .A(N3496), .B(N6952));
NOR2XL inst_cellmath__63_0_I2109 (.Y(N7373), .A(N3702), .B(N6998));
NOR2XL inst_cellmath__63_0_I2091 (.Y(N7345), .A(N3611), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2443 (.CO(N7307), .S(N7116), .A(N7373), .B(N7345), .CI(N3446));
ADDFX1 inst_cellmath__63_0_I2453 (.CO(N7624), .S(N7431), .A(N7022), .B(N6990), .CI(N7307));
NOR2XL inst_cellmath__63_0_I2146 (.Y(N6933), .A(N3432), .B(N7304));
NAND2XL inst_cellmath__63_0_I2218 (.Y(N7051), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[11]));
NOR2XL inst_cellmath__63_0_I2164 (.Y(N6961), .A(N3462), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2452 (.CO(N7236), .S(N7048), .A(N6933), .B(N7051), .CI(N6961));
NOR2XL inst_cellmath__63_0_I2090 (.Y(N6958), .A(N3611), .B(N6998));
NOR2XL inst_cellmath__63_0_I2072 (.Y(N6929), .A(N3446), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2434 (.CO(N7370), .S(N7176), .A(N6958), .B(N6929), .CI(N3412));
NOR2XL inst_cellmath__63_0_I2108 (.Y(N6988), .A(N3702), .B(N7304));
NAND2XL inst_cellmath__63_0_I2216 (.Y(N7160), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[9]));
NOR2XL inst_cellmath__63_0_I2126 (.Y(N7019), .A(N3399), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2435 (.CO(N6871), .S(N7563), .A(N6988), .B(N7160), .CI(N7019));
ADDFX1 inst_cellmath__63_0_I2446 (.CO(N7579), .S(N7383), .A(N7116), .B(N7370), .CI(N6871));
ADDFX1 inst_cellmath__63_0_I2455 (.CO(N7516), .S(N7318), .A(N7431), .B(N7048), .CI(N7579));
ADDFX1 inst_cellmath__63_0_I2462 (.CO(N7560), .S(N7368), .A(N7484), .B(N7128), .CI(N7516));
ADDFX1 inst_cellmath__63_0_I2461 (.CO(N7174), .S(N6981), .A(N7624), .B(N7236), .CI(N7097));
ADDFX1 inst_cellmath__63_0_I2468 (.CO(inst_cellmath__63__W1[29]), .S(inst_cellmath__63__W1[28]), .A(N7560), .B(N7174), .CI(N7530));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1487 (.Y(N4238), .A0(N4533), .A1(N4252), .B0(N4260), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1429 (.Y(N4277), .A0(N4533), .A1(N5159), .B0(N4856), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1535 (.Y(N4415), .A0(N4896), .A1(N4238), .B0(N4277), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I996 (.Y(N4784), .A0(N13807), .A1(N4953), .B0(N13766), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1279 (.Y(N4182), .A0(N4314), .A1(N4869), .B0(N13766), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1323 (.Y(N5111), .A0(N4533), .A1(N4784), .B0(N4182), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1262 (.Y(N4196), .A0(N4533), .A1(N4266), .B0(N5010), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1372 (.Y(N5066), .A0(N4896), .A1(N5111), .B0(N4196), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1587 (.Y(N5080), .A0(N4634), .A1(N4415), .B0(N5066), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1106 (.Y(N4284), .A0(N4533), .A1(N4154), .B0(N4510), .B1(a_man[19]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I986 (.Y(N4202), .A(N4297));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1034 (.Y(N4798), .A0(N4533), .A1(N4915), .B0(N4202), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1152 (.Y(N4460), .A0(N4896), .A1(N4284), .B0(N4798), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I842 (.Y(N4687), .A0(N4280), .A1(N13803), .B0(a_man[17]), .B1(N4826));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I908 (.Y(N4321), .A0(a_man[17]), .A1(N4533), .B0(N4687), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I810 (.Y(N4664), .A0(N4533), .A1(N4958), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I956 (.Y(N4278), .A0(N4896), .A1(N4321), .B0(N4664), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1207 (.Y(N4640), .A0(N4634), .A1(N4460), .B0(N4278), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1640 (.Y(N490), .A0(N4911), .A1(N5080), .B0(N4640), .B1(a_man[22]));
NOR2XL inst_cellmath__63_0_I2198 (.Y(N7136), .A(N3538), .B(N6983));
NOR2XL inst_cellmath__63_0_I2144 (.Y(N7049), .A(N3432), .B(N6952));
NOR2XL inst_cellmath__63_0_I2162 (.Y(N7078), .A(N3462), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2436 (.CO(N7258), .S(N7068), .A(N7136), .B(N7049), .CI(N7078));
NOR2XL inst_cellmath__63_0_I2071 (.Y(N7429), .A(N3446), .B(N6998));
NOR2XL inst_cellmath__63_0_I2053 (.Y(N7399), .A(N3412), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2424 (.CO(N7054), .S(N6856), .A(N7429), .B(N7399), .CI(N3456));
NOR2XL inst_cellmath__63_0_I2180 (.Y(N7107), .A(N3496), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2437 (.CO(N7646), .S(N7454), .A(N7054), .B(N7107), .CI(N7176));
ADDFX1 inst_cellmath__63_0_I2447 (.CO(N7082), .S(N6887), .A(N7502), .B(N7258), .CI(N7646));
ADDFX1 inst_cellmath__63_0_I2456 (.CO(N7013), .S(N7706), .A(N7082), .B(N6932), .CI(N7318));
ADDFX1 inst_cellmath__63_0_I2463 (.CO(inst_cellmath__63__W0[28]), .S(inst_cellmath__63__W1[27]), .A(N7013), .B(N6981), .CI(N7368));
ADDHX1 inst_cellmath__64_0_I2561 (.CO(N8648), .S(N9231), .A(N490), .B(inst_cellmath__63__W0[28]));
ADDFX1 inst_cellmath__64_0_I2566 (.CO(N8773), .S(N8613), .A(N9039), .B(inst_cellmath__63__W1[29]), .CI(N8648));
NAND2XL inst_cellmath__64_0_I2729 (.Y(N8960), .A(N9180), .B(N8773));
NAND2XL inst_cellmath__64_0_I2761 (.Y(N8589), .A(N9273), .B(N8960));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1448 (.Y(N4636), .A0(N4314), .A1(N4166), .B0(N4297), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1486 (.Y(N5036), .A0(N4533), .A1(N4636), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1428 (.Y(N5070), .A0(N4533), .A1(N4172), .B0(N4903), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1534 (.Y(N4193), .A0(N4896), .A1(N5036), .B0(N5070), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1322 (.Y(N4885), .A0(N4533), .A1(N4739), .B0(N4534), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1261 (.Y(N4991), .A0(N4533), .A1(N4457), .B0(N5108), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1371 (.Y(N4841), .A0(N4896), .A1(N4885), .B0(N4991), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1586 (.Y(N4858), .A0(N4634), .A1(N4193), .B0(N4841), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1105 (.Y(N5077), .A0(N4533), .A1(N4357), .B0(N4650), .B1(a_man[19]));
INVXL inst_noninc_a_cellmath__55_2WWMM_I998 (.Y(N5100), .A(N4166));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1033 (.Y(N4571), .A0(N4533), .A1(N5100), .B0(N4998), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1151 (.Y(N4237), .A0(N4896), .A1(N5077), .B0(N4571), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I907 (.Y(N5118), .A0(N4533), .A1(N4929), .B0(N4967), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I809 (.Y(N4441), .A0(N4533), .A1(N4510), .B0(N4717), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I955 (.Y(N5071), .A0(N4896), .A1(N5118), .B0(N4441), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1206 (.Y(N4414), .A0(N4634), .A1(N4237), .B0(N5071), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1639 (.Y(N489), .A0(N4911), .A1(N4858), .B0(N4414), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2557 (.CO(N8830), .S(N8675), .A(N489), .B(inst_cellmath__63__W1[27]));
ADDFX1 inst_cellmath__64_0_I2562 (.CO(N8978), .S(N8802), .A(N9231), .B(inst_cellmath__63__W1[28]), .CI(N8830));
NAND2XL inst_cellmath__64_0_I2727 (.Y(N8630), .A(N8613), .B(N8978));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I870 (.Y(N4877), .A(N13803), .B(N4438));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1484 (.Y(N4591), .A0(N4533), .A1(N4855), .B0(N4877), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1426 (.Y(N4623), .A0(N4875), .A1(N4533), .B0(a_man[19]), .B1(N4805));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1532 (.Y(N4765), .A0(N4896), .A1(N4591), .B0(N4623), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1320 (.Y(N4440), .A0(N4533), .A1(N4918), .B0(N4706), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1259 (.Y(N4544), .A0(N4533), .A1(N4314), .B0(N4981), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1369 (.Y(N4394), .A0(N4896), .A1(N4440), .B0(N4544), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1584 (.Y(N4412), .A0(N4634), .A1(N4765), .B0(N4394), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1068 (.Y(N4937), .A0(N13807), .A1(N4736), .B0(N13764), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1103 (.Y(N4635), .A0(N4533), .A1(N4937), .B0(N4151), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I983 (.Y(N4551), .A0(N13795), .A1(N4280), .B0(N4736), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1031 (.Y(N5152), .A0(N4533), .A1(N4218), .B0(N4551), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1149 (.Y(N4812), .A0(N4896), .A1(N4635), .B0(N5152), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I905 (.Y(N4446), .A0(N4533), .A1(N4877), .B0(N5108), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I807 (.Y(N5013), .A0(N4533), .A1(N4517), .B0(N4739), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I953 (.Y(N4624), .A0(N4896), .A1(N4446), .B0(N5013), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1204 (.Y(N4989), .A0(N4634), .A1(N4812), .B0(N4624), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1637 (.Y(N487), .A0(N4911), .A1(N4412), .B0(N4989), .B1(a_man[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1442 (.Y(N4299), .A(N13772), .B(N4280));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1483 (.Y(N4365), .A0(N4533), .A1(N4652), .B0(N4299), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1392 (.Y(N4573), .A0(N4314), .A1(N4297), .B0(N4869), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1425 (.Y(N4398), .A0(N4533), .A1(N4573), .B0(N5131), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1531 (.Y(N4542), .A0(N4896), .A1(N4365), .B0(N4398), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1319 (.Y(N4215), .A0(N4533), .A1(N4170), .B0(N4188), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1228 (.Y(N5076), .A0(N4314), .A1(a_man[17]), .B0(N4280), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1258 (.Y(N4330), .A0(N4533), .A1(N5076), .B0(N4510), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1368 (.Y(N4173), .A0(N4896), .A1(N4215), .B0(N4330), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1583 (.Y(N4191), .A0(N4634), .A1(N4542), .B0(N4173), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1067 (.Y(N4708), .A0(N13807), .A1(N4300), .B0(N13764), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1102 (.Y(N4410), .A0(N4533), .A1(N4708), .B0(N4377), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1030 (.Y(N4932), .A0(N4533), .A1(N4551), .B0(N4341), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1148 (.Y(N4590), .A0(N4896), .A1(N4410), .B0(N4932), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I904 (.Y(N4224), .A0(N4533), .A1(N4805), .B0(N5108), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I806 (.Y(N4792), .A0(N4533), .A1(N4303), .B0(N4849), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I952 (.Y(N4399), .A0(N4896), .A1(N4224), .B0(N4792), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1203 (.Y(N4764), .A0(N4634), .A1(N4590), .B0(N4399), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1636 (.Y(N486), .A0(N4911), .A1(N4191), .B0(N4764), .B1(a_man[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1482 (.Y(N4148), .A0(N4533), .A1(N5076), .B0(N4584), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1393 (.Y(N4799), .A0(N4314), .A1(N4166), .B0(N4438), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1424 (.Y(N4178), .A0(N4533), .A1(N4799), .B0(N4218), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1530 (.Y(N4328), .A0(N4896), .A1(N4148), .B0(N4178), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1276 (.Y(N4222), .A0(N4314), .A1(N4300), .B0(N4479), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1318 (.Y(N5012), .A0(N4533), .A1(N4572), .B0(N4222), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1257 (.Y(N5129), .A0(N4533), .A1(N4988), .B0(N4188), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1367 (.Y(N4972), .A0(N4896), .A1(N5012), .B0(N5129), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1582 (.Y(N4987), .A0(N4634), .A1(N4328), .B0(N4972), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1101 (.Y(N4187), .A0(N4533), .A1(N4969), .B0(N4958), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I997 (.Y(N5005), .A0(N13807), .A1(N13760), .B0(N4297), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1029 (.Y(N4702), .A0(N4533), .A1(N5005), .B0(N4915), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1147 (.Y(N4364), .A0(N4896), .A1(N4187), .B0(N4702), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I903 (.Y(N5021), .A0(N4533), .A1(N4428), .B0(N4271), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I805 (.Y(N4565), .A0(N4533), .A1(N5061), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I951 (.Y(N4179), .A0(N4896), .A1(N5021), .B0(N4565), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1202 (.Y(N4541), .A0(N4634), .A1(N4364), .B0(N4179), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1635 (.Y(N485), .A0(N4911), .A1(N4987), .B0(N4541), .B1(a_man[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5896 (.Y(N4945), .A0(N4533), .A1(N4573), .B0(N4619), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1423 (.Y(N4977), .A0(N4533), .A1(N4573), .B0(N5101), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5897 (.Y(N5126), .A0(N4896), .A1(N4945), .B0(N4977), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1317 (.Y(N4791), .A0(N4533), .A1(N5140), .B0(N4855), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1256 (.Y(N4902), .A0(N4533), .A1(N4409), .B0(N4971), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1366 (.Y(N4746), .A0(N4896), .A1(N4791), .B0(N4902), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5898 (.Y(N4763), .A0(N4634), .A1(N5126), .B0(N4746), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1100 (.Y(N4984), .A0(N4533), .A1(N4270), .B0(N4154), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I982 (.Y(N4465), .A0(N13795), .A1(N4953), .B0(N4166), .B1(N13782));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1028 (.Y(N4486), .A0(N4533), .A1(N4784), .B0(N4465), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1146 (.Y(N4147), .A0(N4896), .A1(N4984), .B0(N4486), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I902 (.Y(N4800), .A0(N4533), .A1(N4561), .B0(N4531), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I804 (.Y(N4347), .A0(N4533), .A1(N4981), .B0(N4535), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I950 (.Y(N4978), .A0(N4896), .A1(N4800), .B0(N4347), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1201 (.Y(N4327), .A0(N4634), .A1(N4147), .B0(N4978), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I5900 (.Y(N484), .A0(N4911), .A1(N4763), .B0(N4327), .B1(a_man[22]));
ADDHX1 inst_cellmath__64_0_I2535 (.CO(N9142), .S(N8980), .A(N484), .B(N8574));
ADDHX1 inst_cellmath__64_0_I2539 (.CO(N8953), .S(N8777), .A(N485), .B(N9142));
ADDHX1 inst_cellmath__64_0_I2543 (.CO(N8754), .S(N8586), .A(N486), .B(N8953));
ADDHX1 inst_cellmath__64_0_I2548 (.CO(N8893), .S(N8731), .A(N487), .B(N8754));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1485 (.Y(N4813), .A0(N4533), .A1(N5078), .B0(N4903), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1427 (.Y(N4845), .A0(N4533), .A1(N4409), .B0(N4402), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1533 (.Y(N4990), .A0(N4896), .A1(N4813), .B0(N4845), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1277 (.Y(N4318), .A0(N4314), .A1(N4300), .B0(N4166), .B1(N13786));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1321 (.Y(N4663), .A0(N4533), .A1(N4271), .B0(N4318), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1260 (.Y(N4767), .A0(N4533), .A1(N4616), .B0(N4177), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1370 (.Y(N4618), .A0(N4896), .A1(N4663), .B0(N4767), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1585 (.Y(N4639), .A0(N4634), .A1(N4990), .B0(N4618), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1104 (.Y(N4854), .A0(N4533), .A1(N4471), .B0(N4469), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1032 (.Y(N4352), .A0(N4533), .A1(N4341), .B0(N4774), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1150 (.Y(N5035), .A0(N4896), .A1(N4854), .B0(N4352), .B1(a_man[20]));
NAND2BXL inst_noninc_a_cellmath__55_2WWMM_I906 (.Y(N4671), .AN(N4900), .B(N4533));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I808 (.Y(N4216), .A0(N4533), .A1(N4740), .B0(N4501), .B1(a_man[19]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I954 (.Y(N4846), .A0(N4896), .A1(N4671), .B0(N4216), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1205 (.Y(N4192), .A0(N4634), .A1(N5035), .B0(N4846), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1638 (.Y(N488), .A0(N4911), .A1(N4639), .B0(N4192), .B1(a_man[22]));
NOR2XL inst_cellmath__63_0_I2070 (.Y(N7046), .A(N3446), .B(N7304));
NAND2XL inst_cellmath__63_0_I2214 (.Y(N7271), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[7]));
NOR2XL inst_cellmath__63_0_I2196 (.Y(N7244), .A(N3538), .B(N7594));
ADDFX1 inst_cellmath__63_0_I2414 (.CO(N7616), .S(N7422), .A(N7046), .B(N7271), .CI(N7244));
NOR2XL inst_cellmath__63_0_I2106 (.Y(N7105), .A(N3702), .B(N6952));
NOR2XL inst_cellmath__63_0_I2088 (.Y(N7075), .A(N3611), .B(N7533));
NOR2XL inst_cellmath__63_0_I2124 (.Y(N7133), .A(N3399), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2415 (.CO(N7121), .S(N6923), .A(N7105), .B(N7075), .CI(N7133));
ADDFX1 inst_cellmath__63_0_I2428 (.CO(N7712), .S(N7519), .A(N7616), .B(N6856), .CI(N7121));
ADDFX1 inst_cellmath__63_0_I2439 (.CO(N7535), .S(N7340), .A(N7068), .B(N7563), .CI(N7712));
NOR2XL inst_cellmath__63_0_I2052 (.Y(N7014), .A(N3412), .B(N6998));
NOR2XL inst_cellmath__63_0_I2034 (.Y(N6986), .A(N3456), .B(N7576));
ADDFX1 inst_cellmath__63_0_I2413 (.CO(N7227), .S(N7039), .A(N7014), .B(N6986), .CI(N3503));
ADDFX1 inst_cellmath__63_0_I2417 (.CO(N7005), .S(N7697), .A(N7039), .B(N7023), .CI(N7407));
NOR2XL inst_cellmath__63_0_I2161 (.Y(N7574), .A(N3462), .B(N7562));
NOR2XL inst_cellmath__63_0_I2143 (.Y(N7545), .A(N3432), .B(N7257));
ADDFX1 inst_cellmath__63_0_I2427 (.CO(N7325), .S(N7132), .A(N7574), .B(N7545), .CI(N7227));
ADDFX1 inst_cellmath__63_0_I2418 (.CO(N7388), .S(N7196), .A(N7294), .B(N6910), .CI(N7422));
ADDFX1 inst_cellmath__63_0_I2430 (.CO(N7598), .S(N7401), .A(N7005), .B(N7132), .CI(N7388));
NOR2XL inst_cellmath__63_0_I2160 (.Y(N7189), .A(N3462), .B(N6983));
NOR2XL inst_cellmath__63_0_I2178 (.Y(N7216), .A(N3496), .B(N7288));
NOR2XL inst_cellmath__63_0_I2142 (.Y(N7157), .A(N3432), .B(N7562));
ADDFX1 inst_cellmath__63_0_I2416 (.CO(N7507), .S(N7311), .A(N7189), .B(N7216), .CI(N7157));
ADDFX1 inst_cellmath__63_0_I2419 (.CO(N6893), .S(N7582), .A(N7311), .B(N6923), .CI(N7682));
NOR2XL inst_cellmath__63_0_I2089 (.Y(N7460), .A(N3611), .B(N7304));
NAND2XL inst_cellmath__63_0_I2215 (.Y(N7664), .A(inst_cellmath__48[15]), .B(inst_cellmath__51[8]));
NOR2XL inst_cellmath__63_0_I2107 (.Y(N7489), .A(N3702), .B(N7533));
ADDFX1 inst_cellmath__63_0_I2425 (.CO(N7437), .S(N7240), .A(N7460), .B(N7664), .CI(N7489));
NOR2XL inst_cellmath__63_0_I2197 (.Y(N7633), .A(N3538), .B(N7288));
NOR2XL inst_cellmath__63_0_I2125 (.Y(N7520), .A(N3399), .B(N6952));
NOR2XL inst_cellmath__63_0_I2179 (.Y(N7604), .A(N3496), .B(N6983));
ADDFX1 inst_cellmath__63_0_I2426 (.CO(N6937), .S(N7629), .A(N7633), .B(N7520), .CI(N7604));
ADDFX1 inst_cellmath__63_0_I2429 (.CO(N7208), .S(N7018), .A(N7507), .B(N7240), .CI(N7629));
ADDFX1 inst_cellmath__63_0_I2431 (.CO(N7101), .S(N6904), .A(N6893), .B(N7519), .CI(N7018));
ADDFX1 inst_cellmath__63_0_I2441 (.CO(N7419), .S(N7223), .A(N7340), .B(N7598), .CI(N7101));
ADDFX1 inst_cellmath__63_0_I2438 (.CO(N7149), .S(N6953), .A(N6937), .B(N7437), .CI(N7325));
ADDFX1 inst_cellmath__63_0_I2448 (.CO(N7468), .S(N7268), .A(N7149), .B(N7000), .CI(N7383));
ADDFX1 inst_cellmath__63_0_I2440 (.CO(N7035), .S(N6843), .A(N7208), .B(N7454), .CI(N6953));
ADDFX1 inst_cellmath__63_0_I2449 (.CO(N6964), .S(N7660), .A(N6887), .B(N7535), .CI(N7035));
ADDFX1 inst_cellmath__63_0_I2450 (.CO(inst_cellmath__63__W0[26]), .S(inst_cellmath__63__W1[25]), .A(N7419), .B(N7268), .CI(N7660));
ADDFX1 inst_cellmath__64_0_I2553 (.CO(N9029), .S(N8862), .A(N8893), .B(N488), .CI(inst_cellmath__63__W0[26]));
ADDFX1 inst_cellmath__63_0_I2457 (.CO(inst_cellmath__63__W0[27]), .S(inst_cellmath__63__W1[26]), .A(N6964), .B(N7468), .CI(N7706));
ADDFX1 inst_cellmath__64_0_I2558 (.CO(N9168), .S(N9003), .A(N9029), .B(inst_cellmath__63__W0[27]), .CI(N8675));
NAND2XL inst_cellmath__64_0_I2725 (.Y(N9047), .A(N8802), .B(N9168));
NAND2XL inst_cellmath__64_0_I2758 (.Y(N8695), .A(N8630), .B(N9047));
NOR2XL inst_cellmath__64_0_I2763 (.Y(N9156), .A(N8589), .B(N8695));
NAND2XL inst_cellmath__64_0_I2796 (.Y(N9030), .A(N8768), .B(N9156));
NOR2XL inst_cellmath__62_0_I1794 (.Y(inst_cellmath__62__W0[24]), .A(N6347), .B(N6286));
NOR2XL inst_cellmath__62_0_I1793 (.Y(N6329), .A(N6347), .B(N6213));
NOR2XL inst_cellmath__62_0_I1781 (.Y(N6264), .A(N6276), .B(N6286));
NOR2XL inst_cellmath__62_0_I1792 (.Y(N6182), .A(N6347), .B(N6477));
NOR2XL inst_cellmath__62_0_I1768 (.Y(N6385), .A(N6198), .B(N6286));
NOR2XL inst_cellmath__62_0_I1780 (.Y(N6451), .A(N6276), .B(N6213));
ADDFX1 inst_cellmath__62_0_I1880 (.CO(N6459), .S(N6383), .A(N6182), .B(N6385), .CI(N6451));
ADDFX1 inst_cellmath__62_0_I1882 (.CO(inst_cellmath__62__W1[24]), .S(inst_cellmath__62__W0[23]), .A(N6329), .B(N6264), .CI(N6459));
ADDFX1 inst_cellmath__64_0_I2544 (.CO(N9081), .S(N8925), .A(inst_cellmath__62__W0[24]), .B(N8586), .CI(inst_cellmath__62__W1[24]));
ADDFX1 inst_cellmath__63_0_I2420 (.CO(N7274), .S(N7087), .A(N7697), .B(N7181), .CI(N7566));
ADDFX1 inst_cellmath__63_0_I2421 (.CO(N7666), .S(N7472), .A(N7071), .B(N7196), .CI(N7582));
ADDFX1 inst_cellmath__63_0_I2432 (.CO(N7486), .S(N7289), .A(N7401), .B(N7274), .CI(N7666));
ADDFX1 inst_cellmath__63_0_I2442 (.CO(inst_cellmath__63__W0[25]), .S(inst_cellmath__63__W1[24]), .A(N6843), .B(N7486), .CI(N7223));
ADDFX1 inst_cellmath__64_0_I2549 (.CO(N9221), .S(N9054), .A(N9081), .B(N8731), .CI(inst_cellmath__63__W0[25]));
ADDFX1 inst_cellmath__64_0_I2554 (.CO(N8600), .S(N9193), .A(N9221), .B(inst_cellmath__63__W1[26]), .CI(N8862));
NAND2XL inst_cellmath__64_0_I2723 (.Y(N8724), .A(N8600), .B(N9003));
ADDFX1 inst_cellmath__63_0_I2422 (.CO(N7162), .S(N6968), .A(N7087), .B(N7456), .CI(N6955));
ADDFX1 inst_cellmath__63_0_I2433 (.CO(inst_cellmath__63__W0[24]), .S(inst_cellmath__63__W1[23]), .A(N7162), .B(N6904), .CI(N7289));
ADDFX1 inst_cellmath__64_0_I2545 (.CO(N8664), .S(N9244), .A(N8925), .B(inst_cellmath__63__W0[24]), .CI(inst_cellmath__63__W1[24]));
ADDFX1 inst_cellmath__64_0_I2550 (.CO(N8790), .S(N8634), .A(N9054), .B(inst_cellmath__63__W1[25]), .CI(N8664));
NAND2XL inst_cellmath__64_0_I2721 (.Y(N9150), .A(N8790), .B(N9193));
NAND2X1 inst_cellmath__64_0_I2754 (.Y(N8983), .A(N8724), .B(N9150));
ADDFXL inst_cellmath__62_0_I1881 (.CO(inst_cellmath__62__W1[23]), .S(inst_cellmath__62__W0[22]), .A(N6383), .B(N6355), .CI(N6502));
ADDFX1 inst_cellmath__64_0_I2540 (.CO(N9267), .S(N9110), .A(inst_cellmath__62__W0[23]), .B(N8777), .CI(inst_cellmath__62__W1[23]));
ADDFX1 inst_cellmath__63_0_I2423 (.CO(inst_cellmath__63__W0[23]), .S(inst_cellmath__63__W1[22]), .A(N7342), .B(N7472), .CI(N6968));
ADDFX1 inst_cellmath__64_0_I2541 (.CO(N8848), .S(N8690), .A(inst_cellmath__63__W0[23]), .B(inst_cellmath__63__W1[23]), .CI(N9110));
ADDFX1 inst_cellmath__64_0_I2546 (.CO(N8991), .S(N8818), .A(N9267), .B(N9244), .CI(N8848));
NAND2XL inst_cellmath__64_0_I2719 (.Y(N8811), .A(N8634), .B(N8991));
ADDFHXL inst_cellmath__64_0_I2536 (.CO(N8718), .S(N9294), .A(N8980), .B(inst_cellmath__62__W0[22]), .CI(inst_cellmath__63__W0[22]));
ADDFHXL inst_cellmath__64_0_I2537 (.CO(N9042), .S(N8881), .A(inst_cellmath__63__W1[22]), .B(inst_cellmath__62__W1[22]), .CI(N9294));
ADDFX1 inst_cellmath__64_0_I2542 (.CO(N9182), .S(N9017), .A(N8690), .B(N8718), .CI(N9042));
NAND2X1 inst_cellmath__64_0_I2717 (.Y(N9239), .A(N8818), .B(N9182));
NAND2X1 inst_cellmath__64_0_I2751 (.Y(N9071), .A(N8811), .B(N9239));
NOR2X2 inst_cellmath__64_0_I2756 (.Y(N8778), .A(N8983), .B(N9071));
ADDFHXL inst_cellmath__64_0_I2538 (.CO(N8619), .S(N9209), .A(N8913), .B(N9235), .CI(N8881));
NAND2X2 inst_cellmath__64_0_I2715 (.Y(N8922), .A(N8619), .B(N9017));
NOR2X2 inst_cellmath__64_0_I2712 (.Y(N9179), .A(N8805), .B(N9209));
NOR2XL inst_cellmath__64_0_I2714 (.Y(N8750), .A(N8619), .B(N9017));
AOI21X2 inst_cellmath__64_0_I2749 (.Y(N9010), .A0(N8922), .A1(N9179), .B0(N8750));
INVX2 inst_cellmath__64_0_I2781 (.Y(N8828), .A(N9010));
NOR2X1 inst_cellmath__64_0_I2716 (.Y(N9075), .A(N8818), .B(N9182));
NOR2XL inst_cellmath__64_0_I2718 (.Y(N8661), .A(N8634), .B(N8991));
AOI21X2 inst_cellmath__64_0_I2750 (.Y(N8917), .A0(N8811), .A1(N9075), .B0(N8661));
NOR2XL inst_cellmath__64_0_I2720 (.Y(N8986), .A(N8790), .B(N9193));
NOR2XL inst_cellmath__64_0_I2722 (.Y(N9299), .A(N8600), .B(N9003));
AOI21XL inst_cellmath__64_0_I2753 (.Y(N8806), .A0(N8724), .A1(N8986), .B0(N9299));
OAI21X1 inst_cellmath__64_0_I2755 (.Y(N8622), .A0(N8983), .A1(N8917), .B0(N8806));
AOI21X4 inst_cellmath__64_0_I2791 (.Y(N8964), .A0(N8778), .A1(N8828), .B0(N8622));
NOR2XL inst_cellmath__64_0_I2724 (.Y(N8889), .A(N8802), .B(N9168));
NOR2XL inst_cellmath__64_0_I2726 (.Y(N9214), .A(N8613), .B(N8978));
AOI21XL inst_cellmath__64_0_I2757 (.Y(N9268), .A0(N8630), .A1(N8889), .B0(N9214));
NOR2XL inst_cellmath__64_0_I2728 (.Y(N8783), .A(N9180), .B(N8773));
NOR2XL inst_cellmath__64_0_I2730 (.Y(N9120), .A(N8988), .B(N8581));
AOI21XL inst_cellmath__64_0_I2760 (.Y(N9185), .A0(N9273), .A1(N8783), .B0(N9120));
OAI21XL inst_cellmath__64_0_I2762 (.Y(N8993), .A0(N8589), .A1(N9268), .B0(N9185));
NOR2XL inst_cellmath__64_0_I16082 (.Y(N8698), .A(N26158), .B(N26147));
NOR2XL inst_cellmath__64_0_I2734 (.Y(N9023), .A(N8597), .B(N8963));
AOI21XL inst_cellmath__64_0_I2764 (.Y(N8897), .A0(N9189), .A1(N8698), .B0(N9023));
NOR2XL inst_cellmath__64_0_I2736 (.Y(N8596), .A(N9164), .B(N8764));
NOR2XL inst_cellmath__64_0_I2738 (.Y(N8933), .A(N8976), .B(N8567));
AOI21XL inst_cellmath__64_0_I2767 (.Y(N8793), .A0(N9090), .A1(N8596), .B0(N8933));
OAI21XL inst_cellmath__64_0_I2769 (.Y(N8604), .A0(N8969), .A1(N8897), .B0(N8793));
AOI21XL inst_cellmath__64_0_I2795 (.Y(N8861), .A0(N8768), .A1(N8993), .B0(N8604));
OAI21X2 cynw_cm_float_rcp_I16260 (.Y(N26703), .A0(N9030), .A1(N8964), .B0(N8861));
NAND2X2 inst_cellmath__64_0_I2713 (.Y(N8578), .A(N8805), .B(N9209));
CLKAND2X3 inst_cellmath__64_0_I2782 (.Y(N8568), .A(N8922), .B(N8578));
NAND2X2 inst_cellmath__64_0_I2792 (.Y(N9125), .A(N8778), .B(N8568));
NOR2X1 cynw_cm_float_rcp_I16261 (.Y(N26710), .A(N9030), .B(N9125));
AOI21X4 cynw_cm_float_rcp_I16262 (.Y(N8842), .A0(N26710), .A1(N8674), .B0(N26703));
NAND2BXL cynw_cm_float_rcp_I16263 (.Y(N26692), .AN(N9251), .B(N8670));
XOR2XL cynw_cm_float_rcp_I16264 (.Y(N26698), .A(N26692), .B(N8842));
INVXL cynw_cm_float_rcp_I16265 (.Y(N9934), .A(inst_cellmath__67));
AOI22XL cynw_cm_float_rcp_I16266 (.Y(x[19]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(N26698));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I965 (.Y(N4232), .A(a_man[20]), .B(N4718));
OAI2BB1X1 inst_noninc_a_cellmath__55_2WWMM_I1161 (.Y(N4418), .A0N(N5163), .A1N(a_man[19]), .B0(N4896));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1216 (.Y(N4600), .A0(N4634), .A1(N4418), .B0(N4232), .B1(a_man[21]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1217 (.Y(N4821), .A(N4634), .B(N4864));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1270 (.Y(N4824), .A(N4533), .B(N4849));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1381 (.Y(N5025), .A0(N4896), .A1(N4468), .B0(N4824), .B1(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1437 (.Y(N4231), .A0(N4533), .A1(N4341), .B0(N5141), .B1(a_man[19]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1496 (.Y(N4646), .A(N4533), .B(N4968));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1544 (.Y(N4374), .A0(N4896), .A1(N4646), .B0(N4231), .B1(a_man[20]));
NAND2XL inst_noninc_a_cellmath__55_2WWMM_I1545 (.Y(N4601), .A(N4261), .B(a_man[20]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1596 (.Y(N5042), .A0(N4634), .A1(N4374), .B0(N5025), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1597 (.Y(N4246), .A0(N4634), .A1(N4601), .B0(N5093), .B1(a_man[21]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1649 (.Y(N499), .A0(N4911), .A1(N5042), .B0(N4600), .B1(a_man[22]));
AOI22XL inst_noninc_a_cellmath__55_2WWMM_I1650 (.Y(N500), .A0(N4911), .A1(N4246), .B0(N4821), .B1(a_man[22]));
NOR2XL inst_noninc_a_cellmath__55_2WWMM_I1651 (.Y(N4979), .A(N4634), .B(N4964));
OR2XL inst_noninc_a_cellmath__55_2WWMM_I1652 (.Y(N501), .A(N4979), .B(a_man[22]));
OR2XL hap1_A_I6068 (.Y(N8948), .A(1'B0), .B(N498));
INVXL hap1_A_I16319 (.Y(N8576), .A(N499));
OR2XL hap1_A_I6070 (.Y(N8749), .A(1'B0), .B(N499));
INVXL inst_cellmath__64_0_I16320 (.Y(N9147), .A(N500));
NOR2XL inst_cellmath__64_0_I2742 (.Y(N8826), .A(N8948), .B(N8576));
NAND2XL inst_cellmath__64_0_I2743 (.Y(N8998), .A(N8948), .B(N8576));
NOR2XL inst_cellmath__64_0_I2744 (.Y(N9161), .A(N8749), .B(N9147));
NAND2XL inst_cellmath__64_0_I2745 (.Y(N8566), .A(N8749), .B(N9147));
INVXL inst_cellmath__64_0_I2752 (.Y(N9065), .A(N9150));
INVXL inst_cellmath__64_0_I2759 (.Y(N8877), .A(N8960));
INVXL inst_cellmath__64_0_I2766 (.Y(N8688), .A(N8759));
AOI21XL inst_cellmath__64_0_I2771 (.Y(N9258), .A0(N8998), .A1(N9251), .B0(N8826));
NAND2XL inst_cellmath__64_0_I2772 (.Y(N8679), .A(N8998), .B(N8670));
INVXL inst_cellmath__64_0_I2773 (.Y(N9240), .A(N8566));
INVX1 inst_cellmath__64_0_I16084 (.Y(N8741), .A(N8727));
INVXL inst_cellmath__64_0_I2797 (.Y(N8903), .A(N8741));
INVX1 inst_cellmath__64_0_I2798 (.Y(N9064), .A(N9154));
NAND2X2 inst_cellmath__64_0_I16088 (.Y(N8789), .A(N8568), .B(N9092));
AOI21X4 inst_cellmath__64_0_I16085 (.Y(N8730), .A0(N8859), .A1(N9217), .B0(N9122));
AOI21X4 inst_cellmath__64_0_I16087 (.Y(N8635), .A0(N8568), .A1(N8598), .B0(N8828));
OAI21X2 inst_cellmath__64_0_I2801 (.Y(N9004), .A0(N8789), .A1(N8730), .B0(N8635));
NAND2X2 inst_cellmath__64_0_I16086 (.Y(N8894), .A(N8859), .B(N8632));
NOR2X1 inst_cellmath__64_0_I2802 (.Y(N9167), .A(N8789), .B(N8894));
OAI21X2 inst_cellmath__64_0_I2803 (.Y(N8570), .A0(N9125), .A1(N9053), .B0(N8964));
NOR2X1 inst_cellmath__64_0_I2804 (.Y(N8743), .A(N9125), .B(N9220));
INVX1 buf1_A_I6073 (.Y(N13851), .A(N9064));
INVX1 buf1_A_I6074 (.Y(N8643), .A(N13851));
AOI21X2 inst_cellmath__64_0_I2813 (.Y(N8612), .A0(N8903), .A1(N9167), .B0(N9004));
AOI21X2 inst_cellmath__64_0_I2814 (.Y(N8951), .A0(N8743), .A1(N9064), .B0(N8570));
NOR2XL inst_cellmath__64_0_I2817 (.Y(N8696), .A(N9065), .B(N8917));
NOR2XL inst_cellmath__64_0_I2818 (.Y(N9011), .A(N8696), .B(N8986));
NOR2XL inst_cellmath__64_0_I2819 (.Y(N9086), .A(N8877), .B(N9268));
NOR2XL inst_cellmath__64_0_I2820 (.Y(N9237), .A(N9086), .B(N8783));
NOR2XL inst_cellmath__64_0_I2821 (.Y(N8736), .A(N8688), .B(N8897));
NOR2XL inst_cellmath__64_0_I2822 (.Y(N8721), .A(N8736), .B(N8596));
NOR2XL inst_cellmath__64_0_I2823 (.Y(N9129), .A(N9240), .B(N9258));
NOR2XL inst_cellmath__64_0_I2824 (.Y(N8957), .A(N9129), .B(N9161));
NAND2BXL inst_cellmath__64_0_I2827 (.Y(N9117), .AN(N9038), .B(N9206));
NAND2BXL inst_cellmath__64_0_I2828 (.Y(N8854), .AN(N8610), .B(N8772));
NAND2BXL inst_cellmath__64_0_I2829 (.Y(N8592), .AN(N8949), .B(N9103));
NAND2BXL inst_cellmath__64_0_I2830 (.Y(N9087), .AN(N9262), .B(N8686));
NAND2BXL inst_cellmath__64_0_I2831 (.Y(N8823), .AN(N8839), .B(N9013));
NAND2BXL inst_cellmath__64_0_I2832 (.Y(N8563), .AN(N9179), .B(N8578));
NAND2BXL inst_cellmath__64_0_I2833 (.Y(N9060), .AN(N8750), .B(N8922));
NAND2BXL inst_cellmath__64_0_I2834 (.Y(N8796), .AN(N9075), .B(N9239));
NAND2BXL inst_cellmath__64_0_I2835 (.Y(N9284), .AN(N8661), .B(N8811));
NAND2BXL inst_cellmath__64_0_I2836 (.Y(N8956), .AN(N8986), .B(N9150));
NAND2BXL inst_cellmath__64_0_I2837 (.Y(N9247), .AN(N9299), .B(N8724));
NAND2BXL inst_cellmath__64_0_I2838 (.Y(N9259), .AN(N8889), .B(N9047));
NAND2BXL inst_cellmath__64_0_I2839 (.Y(N9008), .AN(N9214), .B(N8630));
NAND2BXL inst_cellmath__64_0_I2840 (.Y(N9198), .AN(N8783), .B(N8960));
NAND2BXL inst_cellmath__64_0_I2841 (.Y(N8746), .AN(N9120), .B(N9273));
NAND2BXL inst_cellmath__64_0_I2843 (.Y(N8719), .AN(N9023), .B(N9189));
NAND2BXL inst_cellmath__64_0_I2844 (.Y(N8691), .AN(N8596), .B(N8759));
NAND2BXL inst_cellmath__64_0_I2845 (.Y(N8992), .AN(N8933), .B(N9090));
NAND2BXL inst_cellmath__64_0_I2847 (.Y(N9183), .AN(N8826), .B(N8998));
NAND2BXL inst_cellmath__64_0_I2848 (.Y(N8939), .AN(N9161), .B(N8566));
XNOR2X1 inst_cellmath__64_0_I16321 (.Y(N9234), .A(N500), .B(N501));
XNOR2X1 inst_cellmath__64_0_I2852 (.Y(inst_cellmath__64[18]), .A(N8854), .B(N8643));
OAI21X4 inst_cellmath__64_0_I16091 (.Y(N9094), .A0(N8894), .A1(N8741), .B0(N8730));
XNOR2X1 inst_cellmath__64_0_I2853 (.Y(inst_cellmath__64[20]), .A(N9094), .B(N9087));
XNOR2X1 inst_cellmath__64_0_I2854 (.Y(inst_cellmath__64[22]), .A(N8674), .B(N8563));
XOR2XL inst_cellmath__64_0_I2855 (.Y(inst_cellmath__64[24]), .A(N8796), .B(N8612));
XOR2XL inst_cellmath__64_0_I2856 (.Y(inst_cellmath__64[28]), .A(N9259), .B(N8951));
AOI21X1 inst_cellmath__64_0_I16089 (.Y(N26156), .A0(N9156), .A1(N8622), .B0(N8993));
NAND2X1 inst_cellmath__64_0_I16090 (.Y(N26165), .A(N9156), .B(N8778));
NOR2X1 inst_cellmath__64_0_I16092 (.Y(N26143), .A(N26165), .B(N8635));
NOR2BX1 inst_cellmath__64_0_I16322 (.Y(N26168), .AN(N26156), .B(N26143));
OAI21X1 inst_cellmath__64_0_I16095 (.Y(N26140), .A0(N26165), .A1(N8635), .B0(N26156));
NOR2X1 inst_cellmath__64_0_I16096 (.Y(N26151), .A(N26165), .B(N8789));
AOI21X2 inst_cellmath__64_0_I16098 (.Y(N9263), .A0(N26151), .A1(N9094), .B0(N26140));
NAND2BXL inst_cellmath__64_0_I16099 (.Y(N26170), .AN(N8698), .B(N8857));
OAI2BB1X1 inst_cellmath__64_0_I16324 (.Y(N26149), .A0N(N26151), .A1N(N9094), .B0(N26168));
INVXL xnor2_A_I16396 (.Y(N26737), .A(N26170));
MXI2XL xnor2_A_I16397 (.Y(inst_cellmath__64[32]), .A(N26170), .B(N26737), .S0(N26149));
XNOR2X1 inst_cellmath__64_0_I2859 (.Y(N9126), .A(N8873), .B(N9117));
XNOR2X1 inst_cellmath__64_0_I2860 (.Y(N8967), .A(N8715), .B(N9117));
MX2XL inst_cellmath__64_0_I2861 (.Y(inst_cellmath__64[17]), .A(N8967), .B(N9126), .S0(N8903));
XNOR2X1 inst_cellmath__64_0_I2862 (.Y(N8863), .A(N8772), .B(N8592));
XNOR2X1 inst_cellmath__64_0_I2863 (.Y(N8705), .A(N8610), .B(N8592));
MX2XL inst_cellmath__64_0_I2864 (.Y(inst_cellmath__64[19]), .A(N8705), .B(N8863), .S0(N8643));
XNOR2X1 inst_cellmath__64_0_I2865 (.Y(N8602), .A(N8686), .B(N8823));
XNOR2X1 inst_cellmath__64_0_I2866 (.Y(N9195), .A(N8823), .B(N9262));
MX2XL inst_cellmath__64_0_I2867 (.Y(inst_cellmath__64[21]), .A(N9195), .B(N8602), .S0(N9094));
XNOR2X1 inst_cellmath__64_0_I2868 (.Y(N9096), .A(N9060), .B(N8578));
XNOR2X1 inst_cellmath__64_0_I2869 (.Y(N8940), .A(N9060), .B(N9179));
MX2XL inst_cellmath__64_0_I2870 (.Y(inst_cellmath__64[23]), .A(N8940), .B(N9096), .S0(N8674));
XNOR2X1 inst_cellmath__64_0_I2871 (.Y(N8831), .A(N9284), .B(N9239));
XNOR2X1 inst_cellmath__64_0_I2872 (.Y(N8677), .A(N9284), .B(N9075));
MX2XL inst_cellmath__64_0_I2873 (.Y(inst_cellmath__64[25]), .A(N8831), .B(N8677), .S0(N8612));
XOR2XL inst_cellmath__64_0_I2874 (.Y(N9170), .A(N8956), .B(N8917));
NAND2XL inst_cellmath__64_0_I2875 (.Y(N8625), .A(N9071), .B(N8917));
XNOR2X1 inst_cellmath__64_0_I2876 (.Y(N8572), .A(N8956), .B(N8625));
MX2XL inst_cellmath__64_0_I2877 (.Y(inst_cellmath__64[26]), .A(N8572), .B(N9170), .S0(N8612));
XOR2XL inst_cellmath__64_0_I2878 (.Y(N8911), .A(N9247), .B(N9011));
OAI21XL inst_cellmath__64_0_I2879 (.Y(N8929), .A0(N9065), .A1(N9071), .B0(N9011));
XNOR2X1 inst_cellmath__64_0_I2880 (.Y(N9068), .A(N9247), .B(N8929));
MX2XL inst_cellmath__64_0_I2881 (.Y(inst_cellmath__64[27]), .A(N9068), .B(N8911), .S0(N8612));
XNOR2X1 inst_cellmath__64_0_I2882 (.Y(N8803), .A(N9008), .B(N9047));
XNOR2X1 inst_cellmath__64_0_I2883 (.Y(N8651), .A(N9008), .B(N8889));
MX2XL inst_cellmath__64_0_I2884 (.Y(inst_cellmath__64[29]), .A(N8803), .B(N8651), .S0(N8951));
XOR2XL inst_cellmath__64_0_I2885 (.Y(N9140), .A(N9198), .B(N9268));
NAND2XL inst_cellmath__64_0_I2886 (.Y(N8867), .A(N8695), .B(N9268));
XNOR2X1 inst_cellmath__64_0_I2887 (.Y(N9292), .A(N9198), .B(N8867));
MX2XL inst_cellmath__64_0_I2888 (.Y(inst_cellmath__64[30]), .A(N9292), .B(N9140), .S0(N8951));
XOR2XL inst_cellmath__64_0_I2889 (.Y(N8879), .A(N8746), .B(N9237));
OAI21XL inst_cellmath__64_0_I2890 (.Y(N9174), .A0(N8877), .A1(N8695), .B0(N9237));
XNOR2X1 inst_cellmath__64_0_I2891 (.Y(N9040), .A(N8746), .B(N9174));
MX2XL inst_cellmath__64_0_I2892 (.Y(inst_cellmath__64[31]), .A(N9040), .B(N8879), .S0(N8951));
XNOR2X1 inst_cellmath__64_0_I2893 (.Y(N8774), .A(N8719), .B(N8857));
XNOR2X1 inst_cellmath__64_0_I2894 (.Y(N8616), .A(N8719), .B(N8698));
MX2XL inst_cellmath__64_0_I2895 (.Y(inst_cellmath__64[33]), .A(N8774), .B(N8616), .S0(N9263));
XOR2XL inst_cellmath__64_0_I2896 (.Y(N9108), .A(N8691), .B(N8897));
NAND2XL inst_cellmath__64_0_I2897 (.Y(N9112), .A(N9057), .B(N8897));
XNOR2X1 inst_cellmath__64_0_I2898 (.Y(N9265), .A(N8691), .B(N9112));
MX2XL inst_cellmath__64_0_I2899 (.Y(inst_cellmath__64[34]), .A(N9265), .B(N9108), .S0(N9263));
XOR2XL inst_cellmath__64_0_I2900 (.Y(N8846), .A(N8992), .B(N8721));
OAI21XL inst_cellmath__64_0_I2901 (.Y(N8665), .A0(N8688), .A1(N9057), .B0(N8721));
XNOR2X1 inst_cellmath__64_0_I2902 (.Y(N9015), .A(N8992), .B(N8665));
MX2XL inst_cellmath__64_0_I2903 (.Y(inst_cellmath__64[35]), .A(N9015), .B(N8846), .S0(N9263));
XNOR2X1 inst_cellmath__64_0_I2904 (.Y(N8752), .A(N9183), .B(N8670));
XNOR2X1 inst_cellmath__64_0_I2905 (.Y(N8584), .A(N9183), .B(N9251));
MX2XL inst_cellmath__64_0_I2906 (.Y(inst_cellmath__64[37]), .A(N8752), .B(N8584), .S0(N8842));
XOR2XL inst_cellmath__64_0_I2907 (.Y(N9080), .A(N8939), .B(N9258));
NAND2XL inst_cellmath__64_0_I2908 (.Y(N8601), .A(N8679), .B(N9258));
XNOR2X1 inst_cellmath__64_0_I2909 (.Y(N9242), .A(N8939), .B(N8601));
MX2XL inst_cellmath__64_0_I2910 (.Y(inst_cellmath__64[38]), .A(N9242), .B(N9080), .S0(N8842));
XOR2XL inst_cellmath__64_0_I2911 (.Y(N8817), .A(N9234), .B(N8957));
OAI21XL inst_cellmath__64_0_I2912 (.Y(N8909), .A0(N9240), .A1(N8679), .B0(N8957));
XNOR2X1 inst_cellmath__64_0_I2913 (.Y(N8989), .A(N9234), .B(N8909));
MX2XL inst_cellmath__64_0_I2914 (.Y(inst_cellmath__64[39]), .A(N8989), .B(N8817), .S0(N8842));
AOI22XL inst_cellmath__68_0_I2940 (.Y(x[0]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[17]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2941 (.Y(x[1]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[18]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2942 (.Y(x[2]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[19]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2943 (.Y(x[3]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[20]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2944 (.Y(x[4]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[21]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2945 (.Y(x[5]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[22]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2946 (.Y(x[6]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__64[23]), .B1(inst_cellmath__67));
AOI22XL inst_cellmath__68_0_I2947 (.Y(x[7]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(inst_cellmath__64[24]));
AOI22XL inst_cellmath__68_0_I2948 (.Y(x[8]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[25]));
AOI22XL inst_cellmath__68_0_I2949 (.Y(x[9]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[26]));
AOI22XL inst_cellmath__68_0_I2950 (.Y(x[10]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[27]));
AOI22XL inst_cellmath__68_0_I2951 (.Y(x[11]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[28]));
AOI22XL inst_cellmath__68_0_I2952 (.Y(x[12]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(inst_cellmath__64[29]));
AOI22XL inst_cellmath__68_0_I2953 (.Y(x[13]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[30]));
AOI22XL inst_cellmath__68_0_I2954 (.Y(x[14]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[31]));
AOI22XL inst_cellmath__68_0_I2955 (.Y(x[15]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(inst_cellmath__64[32]));
AOI22XL inst_cellmath__68_0_I2956 (.Y(x[16]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(inst_cellmath__64[33]));
AOI22XL inst_cellmath__68_0_I2957 (.Y(x[17]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[34]));
AOI22XL inst_cellmath__68_0_I2958 (.Y(x[18]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[35]));
AOI22XL inst_cellmath__68_0_I2960 (.Y(x[20]), .A0(N9934), .A1(N3320), .B0(inst_cellmath__67), .B1(inst_cellmath__64[37]));
AOI22XL inst_cellmath__68_0_I2961 (.Y(x[21]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[38]));
AOI22XL inst_cellmath__68_0_I2962 (.Y(x[22]), .A0(N3320), .A1(N9934), .B0(inst_cellmath__67), .B1(inst_cellmath__64[39]));
assign inst_cellmath__19[1] = 1'B1;
assign inst_cellmath__19[2] = 1'B1;
assign inst_cellmath__19[3] = 1'B1;
assign inst_cellmath__19[4] = 1'B1;
assign inst_cellmath__19[5] = 1'B1;
assign inst_cellmath__19[6] = 1'B1;
assign inst_cellmath__19[7] = 1'B1;
assign inst_cellmath__19[8] = 1'B1;
assign inst_cellmath__48[0] = a_man[0];
assign inst_cellmath__48[1] = a_man[1];
assign inst_cellmath__48[2] = a_man[2];
assign inst_cellmath__48[3] = a_man[3];
assign inst_cellmath__48[4] = a_man[4];
assign inst_cellmath__48[5] = a_man[5];
assign inst_cellmath__48[6] = a_man[6];
assign inst_cellmath__48[7] = a_man[7];
assign inst_cellmath__48[8] = a_man[8];
assign inst_cellmath__48[9] = a_man[9];
assign inst_cellmath__48[10] = a_man[10];
assign inst_cellmath__48[11] = a_man[11];
assign inst_cellmath__48[12] = a_man[12];
assign inst_cellmath__48[13] = a_man[13];
assign inst_cellmath__48[14] = a_man[14];
assign inst_cellmath__51[13] = 1'B0;
assign inst_cellmath__51[14] = 1'B0;
assign inst_cellmath__51[18] = 1'B1;
assign inst_cellmath__60[0] = 1'B0;
assign inst_cellmath__60[1] = 1'B0;
assign inst_cellmath__60[2] = 1'B0;
assign inst_cellmath__60[3] = 1'B0;
assign inst_cellmath__60[4] = 1'B0;
assign inst_cellmath__60[5] = 1'B0;
assign inst_cellmath__60[6] = 1'B0;
assign inst_cellmath__60[7] = 1'B0;
assign inst_cellmath__60[8] = 1'B0;
assign inst_cellmath__60[9] = 1'B0;
assign inst_cellmath__60[10] = 1'B0;
assign inst_cellmath__60[11] = 1'B0;
assign inst_cellmath__60[12] = 1'B0;
assign inst_cellmath__60[13] = 1'B0;
assign inst_cellmath__60[14] = 1'B0;
assign inst_cellmath__60[15] = 1'B0;
assign inst_cellmath__60[16] = 1'B0;
assign inst_cellmath__60[18] = 1'B0;
assign inst_cellmath__60[19] = 1'B0;
assign inst_cellmath__60[20] = 1'B0;
assign inst_cellmath__60[21] = 1'B0;
assign inst_cellmath__60[22] = 1'B0;
assign inst_cellmath__60[23] = 1'B0;
assign inst_cellmath__60[24] = 1'B0;
assign inst_cellmath__62__W0[0] = 1'B0;
assign inst_cellmath__62__W0[1] = 1'B0;
assign inst_cellmath__62__W0[2] = 1'B0;
assign inst_cellmath__62__W0[3] = 1'B0;
assign inst_cellmath__62__W0[8] = 1'B0;
assign inst_cellmath__62__W0[9] = 1'B0;
assign inst_cellmath__62__W0[10] = 1'B0;
assign inst_cellmath__62__W0[15] = 1'B0;
assign inst_cellmath__62__W0[16] = 1'B0;
assign inst_cellmath__62__W0[17] = 1'B0;
assign inst_cellmath__62__W0[25] = 1'B0;
assign inst_cellmath__62__W0[26] = 1'B0;
assign inst_cellmath__62__W0[27] = 1'B0;
assign inst_cellmath__62__W0[28] = 1'B0;
assign inst_cellmath__62__W0[29] = 1'B0;
assign inst_cellmath__62__W0[30] = 1'B0;
assign inst_cellmath__62__W0[31] = 1'B0;
assign inst_cellmath__62__W0[32] = 1'B0;
assign inst_cellmath__62__W0[33] = 1'B0;
assign inst_cellmath__62__W0[34] = 1'B0;
assign inst_cellmath__62__W0[35] = 1'B0;
assign inst_cellmath__62__W0[36] = 1'B0;
assign inst_cellmath__62__W0[37] = 1'B0;
assign inst_cellmath__62__W0[38] = 1'B0;
assign inst_cellmath__62__W0[39] = 1'B0;
assign inst_cellmath__62__W1[0] = 1'B0;
assign inst_cellmath__62__W1[1] = 1'B0;
assign inst_cellmath__62__W1[2] = 1'B0;
assign inst_cellmath__62__W1[3] = 1'B0;
assign inst_cellmath__62__W1[4] = 1'B0;
assign inst_cellmath__62__W1[9] = 1'B0;
assign inst_cellmath__62__W1[10] = 1'B0;
assign inst_cellmath__62__W1[16] = 1'B0;
assign inst_cellmath__62__W1[17] = 1'B0;
assign inst_cellmath__62__W1[25] = 1'B0;
assign inst_cellmath__62__W1[26] = 1'B0;
assign inst_cellmath__62__W1[27] = 1'B0;
assign inst_cellmath__62__W1[28] = 1'B0;
assign inst_cellmath__62__W1[29] = 1'B0;
assign inst_cellmath__62__W1[30] = 1'B0;
assign inst_cellmath__62__W1[31] = 1'B0;
assign inst_cellmath__62__W1[32] = 1'B0;
assign inst_cellmath__62__W1[33] = 1'B0;
assign inst_cellmath__62__W1[34] = 1'B0;
assign inst_cellmath__62__W1[35] = 1'B0;
assign inst_cellmath__62__W1[36] = 1'B0;
assign inst_cellmath__62__W1[37] = 1'B0;
assign inst_cellmath__62__W1[38] = 1'B0;
assign inst_cellmath__62__W1[39] = 1'B0;
assign inst_cellmath__63__W0[0] = 1'B0;
assign inst_cellmath__63__W0[1] = 1'B0;
assign inst_cellmath__63__W0[8] = 1'B0;
assign inst_cellmath__63__W0[9] = 1'B0;
assign inst_cellmath__63__W0[10] = 1'B0;
assign inst_cellmath__63__W0[16] = 1'B0;
assign inst_cellmath__63__W0[17] = 1'B0;
assign inst_cellmath__63__W0[33] = 1'B0;
assign inst_cellmath__63__W0[34] = 1'B1;
assign inst_cellmath__63__W0[35] = 1'B1;
assign inst_cellmath__63__W0[36] = 1'B1;
assign inst_cellmath__63__W0[37] = 1'B1;
assign inst_cellmath__63__W0[38] = 1'B1;
assign inst_cellmath__63__W0[39] = 1'B1;
assign inst_cellmath__63__W1[0] = 1'B0;
assign inst_cellmath__63__W1[1] = 1'B0;
assign inst_cellmath__63__W1[9] = 1'B0;
assign inst_cellmath__63__W1[10] = 1'B0;
assign inst_cellmath__63__W1[15] = 1'B0;
assign inst_cellmath__63__W1[16] = 1'B0;
assign inst_cellmath__63__W1[17] = 1'B0;
assign inst_cellmath__63__W1[34] = 1'B0;
assign inst_cellmath__63__W1[35] = 1'B0;
assign inst_cellmath__63__W1[36] = 1'B0;
assign inst_cellmath__63__W1[37] = 1'B0;
assign inst_cellmath__63__W1[38] = 1'B0;
assign inst_cellmath__63__W1[39] = 1'B0;
assign inst_cellmath__64[0] = 1'B0;
assign inst_cellmath__64[1] = 1'B0;
assign inst_cellmath__64[2] = 1'B0;
assign inst_cellmath__64[3] = 1'B0;
assign inst_cellmath__64[4] = 1'B0;
assign inst_cellmath__64[5] = 1'B0;
assign inst_cellmath__64[6] = 1'B0;
assign inst_cellmath__64[7] = 1'B0;
assign inst_cellmath__64[8] = 1'B0;
assign inst_cellmath__64[9] = 1'B0;
assign inst_cellmath__64[10] = 1'B0;
assign inst_cellmath__64[11] = 1'B0;
assign inst_cellmath__64[12] = 1'B0;
assign inst_cellmath__64[13] = 1'B0;
assign inst_cellmath__64[14] = 1'B0;
assign inst_cellmath__64[15] = 1'B0;
assign inst_cellmath__64[16] = 1'B0;
assign inst_cellmath__64[36] = 1'B0;
assign x[32] = 1'B0;
assign x[33] = 1'B0;
assign x[34] = 1'B0;
assign x[35] = 1'B0;
assign x[36] = 1'B0;
endmodule

/* CADENCE  ubnxQgzarxw= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



