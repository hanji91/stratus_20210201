/*****************************************************************************
    Verilog Hierarchical Gate Level Netlist
    
    Configured at: 22:38:00 KST (+0900), Thursday 31 December 2020
    Configured on: design1
    Configured by: hanji ()
    
    Created by: CellMath Designer 2019.1.01 
*******************************************************************************/
/*****************************************************************************
    Technology library details
    
    name: slow_vdd1v2
    file name(s):
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/generic.lbf
            /usr/cadence/installs/Stratus/tools.lnx86/cellmath/libs/gencount.lbf
            /usr/cadence/installs/Stratus/share/stratus/techlibs/GPDK045/gsclib045_svt_v4.4/gsclib045/timing/slow_vdd1v2_basicCells.lib
    No wireload model
    op condition: PVT_1P08V_125C
*****************************************************************************/

module fp_add_cynw_cm_float_add2_ieee_E8_M23_4_0 (
	a_sign,
	a_exp,
	a_man,
	b_sign,
	b_exp,
	b_man,
	rm,
	x,
	aclk,
	astall
	); /* architecture "gate_level" */ 
input  a_sign;
input [7:0] a_exp;
input [22:0] a_man;
input  b_sign;
input [7:0] b_exp;
input [22:0] b_man;
input [2:0] rm;
output [31:0] x;
input  aclk;
input  astall;
wire  bdw_enable,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18;
wire [8:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35;
wire [49:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37;
wire [25:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44;
wire [26:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
wire [5:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49;
wire [24:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55;
wire [23:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57;
wire [9:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
wire [22:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66;
wire [7:0] fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68;
wire  fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908,
	fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916;
wire N5123,N5130,N5137,N5144,N5151,N5158,N5165 
	,N5172,N5179,N5186,N5193,N5200,N5207,N5214,N5221 
	,N5228,N5235,N5242,N5249,N5256,N5263,N5270,N5334 
	,N5336,N5572,N5588,N5590,N5614,N5616,N5700,N5705 
	,N5974,N6033,N6055,N6057,N6086,N6093,N6095,N6102 
	,N6138,N6147,N6523,N6777,N6784,N6860,N6930,N6937 
	,N6943,N6945,N6947,N6953,N7046,N7165,N7172,N7303 
	,N7323,N7343,N7350,N7357,N7364,N7371,N7379,N7421 
	,N7608,N7662,N7752,N7768,N7820,N7871,N7873,N7941 
	,N7946,N7955,N7962,N7969,N7976,N7983,N7990,N7997 
	,N8003,N8005,N8011,N8013,N8030,N8038,N8046,N8054 
	,N8062,N8070,N8078,N8086,N8148,N8522,N8527,N8533 
	,N8535,N8544,N9015,N9016,N9073,N9074,N9082,N9086 
	,N9088,N9100,N9101,N9115,N9117,N9121,N9123,N9125 
	,N9127,N9128,N9130,N9132,N9135,N9136,N9144,N9147 
	,N9149,N9151,N9156,N9158,N9161,N9163,N9168,N9172 
	,N9205,N9206,N9208,N9213,N9217,N9236,N9238,N9239 
	,N9261,N9265,N9267,N9269,N9273,N9294,N9298,N9303 
	,N9312,N9314,N9318,N9326,N9347,N9348,N9349,N9354 
	,N9355,N9361,N9373,N9377,N9381,N9385,N9387,N9391 
	,N9395,N9397,N9401,N9407,N9410,N9438,N9441,N9445 
	,N9448,N9459,N9464,N9469,N9474;
reg x_reg_22__retimed_I4614_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4614_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3];
	end
assign N8544 = x_reg_22__retimed_I4614_QOUT;
reg x_reg_22__retimed_I4611_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4611_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827;
	end
assign N8535 = x_reg_22__retimed_I4611_QOUT;
reg x_reg_22__retimed_I4610_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4610_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831;
	end
assign N8533 = x_reg_22__retimed_I4610_QOUT;
reg x_reg_22__retimed_I4608_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4608_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7];
	end
assign N8527 = x_reg_22__retimed_I4608_QOUT;
reg x_reg_22__retimed_I4606_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4606_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4];
	end
assign N8522 = x_reg_22__retimed_I4606_QOUT;
reg x_reg_22__retimed_I4437_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4437_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14];
	end
assign N8148 = x_reg_22__retimed_I4437_QOUT;
reg x_reg_22__retimed_I4406_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4406_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679;
	end
assign N8086 = x_reg_22__retimed_I4406_QOUT;
reg x_reg_22__retimed_I4403_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4403_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609;
	end
assign N8078 = x_reg_22__retimed_I4403_QOUT;
reg x_reg_22__retimed_I4400_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4400_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687;
	end
assign N8070 = x_reg_22__retimed_I4400_QOUT;
reg x_reg_22__retimed_I4397_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4397_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618;
	end
assign N8062 = x_reg_22__retimed_I4397_QOUT;
reg x_reg_22__retimed_I4394_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4394_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695;
	end
assign N8054 = x_reg_22__retimed_I4394_QOUT;
reg x_reg_22__retimed_I4391_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4391_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626;
	end
assign N8046 = x_reg_22__retimed_I4391_QOUT;
reg x_reg_22__retimed_I4388_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4388_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704;
	end
assign N8038 = x_reg_22__retimed_I4388_QOUT;
reg x_reg_22__retimed_I4385_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4385_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257;
	end
assign N8030 = x_reg_22__retimed_I4385_QOUT;
reg x_reg_22__retimed_I4380_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4380_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722;
	end
assign N8013 = x_reg_22__retimed_I4380_QOUT;
reg x_reg_22__retimed_I4379_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4379_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664;
	end
assign N8011 = x_reg_22__retimed_I4379_QOUT;
reg x_reg_22__retimed_I4378_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4378_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636;
	end
assign N8005 = x_reg_22__retimed_I4378_QOUT;
reg x_reg_22__retimed_I4377_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4377_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659;
	end
assign N8003 = x_reg_22__retimed_I4377_QOUT;
reg x_reg_22__retimed_I4376_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4376_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700;
	end
assign N7997 = x_reg_22__retimed_I4376_QOUT;
reg x_reg_22__retimed_I4374_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4374_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620;
	end
assign N7990 = x_reg_22__retimed_I4374_QOUT;
reg x_reg_22__retimed_I4372_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4372_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682;
	end
assign N7983 = x_reg_22__retimed_I4372_QOUT;
reg x_reg_22__retimed_I4370_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4370_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600;
	end
assign N7976 = x_reg_22__retimed_I4370_QOUT;
reg x_reg_22__retimed_I4368_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4368_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665;
	end
assign N7969 = x_reg_22__retimed_I4368_QOUT;
reg x_reg_22__retimed_I4366_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4366_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582;
	end
assign N7962 = x_reg_22__retimed_I4366_QOUT;
reg x_reg_22__retimed_I4364_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4364_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644;
	end
assign N7955 = x_reg_22__retimed_I4364_QOUT;
reg x_reg_22__retimed_I4361_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4361_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25];
	end
assign N7946 = x_reg_22__retimed_I4361_QOUT;
reg x_reg_22__retimed_I4360_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4360_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677;
	end
assign N7941 = x_reg_22__retimed_I4360_QOUT;
reg x_reg_22__retimed_I4337_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4337_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894;
	end
assign N7873 = x_reg_22__retimed_I4337_QOUT;
reg x_reg_22__retimed_I4336_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4336_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914;
	end
assign N7871 = x_reg_22__retimed_I4336_QOUT;
reg x_reg_22__retimed_I4318_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4318_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874;
	end
assign N7820 = x_reg_22__retimed_I4318_QOUT;
reg x_reg_22__retimed_I4300_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4300_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840;
	end
assign N7768 = x_reg_22__retimed_I4300_QOUT;
reg x_reg_22__retimed_I4293_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4293_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863;
	end
assign N7752 = x_reg_22__retimed_I4293_QOUT;
reg x_reg_22__retimed_I4272_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4272_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896;
	end
assign N7662 = x_reg_22__retimed_I4272_QOUT;
reg x_reg_22__retimed_I4263_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4263_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845;
	end
assign N7608 = x_reg_22__retimed_I4263_QOUT;
reg x_reg_22__retimed_I4235_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4235_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486;
	end
assign N7421 = x_reg_22__retimed_I4235_QOUT;
reg x_reg_22__retimed_I4221_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4221_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0];
	end
assign N7379 = x_reg_22__retimed_I4221_QOUT;
reg x_reg_22__retimed_I4218_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4218_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1];
	end
assign N7371 = x_reg_22__retimed_I4218_QOUT;
reg x_reg_22__retimed_I4215_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4215_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2];
	end
assign N7364 = x_reg_22__retimed_I4215_QOUT;
reg x_reg_22__retimed_I4212_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4212_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4];
	end
assign N7357 = x_reg_22__retimed_I4212_QOUT;
reg x_reg_22__retimed_I4209_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4209_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5];
	end
assign N7350 = x_reg_22__retimed_I4209_QOUT;
reg x_reg_22__retimed_I4206_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4206_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6];
	end
assign N7343 = x_reg_22__retimed_I4206_QOUT;
reg x_reg_22__retimed_I4198_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4198_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42;
	end
assign N7323 = x_reg_22__retimed_I4198_QOUT;
reg x_reg_22__retimed_I4191_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4191_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3];
	end
assign N7303 = x_reg_22__retimed_I4191_QOUT;
reg x_reg_22__retimed_I4157_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4157_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8];
	end
assign N7172 = x_reg_22__retimed_I4157_QOUT;
reg x_reg_22__retimed_I4154_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4154_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7];
	end
assign N7165 = x_reg_22__retimed_I4154_QOUT;
reg x_reg_22__retimed_I4108_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4108_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4;
	end
assign N7046 = x_reg_22__retimed_I4108_QOUT;
reg x_reg_22__retimed_I4071_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4071_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43;
	end
assign N6953 = x_reg_22__retimed_I4071_QOUT;
reg x_reg_22__retimed_I4069_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4069_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8;
	end
assign N6947 = x_reg_22__retimed_I4069_QOUT;
reg x_reg_22__retimed_I4068_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4068_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635;
	end
assign N6945 = x_reg_22__retimed_I4068_QOUT;
reg x_reg_22__retimed_I4067_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4067_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634;
	end
assign N6943 = x_reg_22__retimed_I4067_QOUT;
reg x_reg_22__retimed_I4065_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4065_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9];
	end
assign N6937 = x_reg_22__retimed_I4065_QOUT;
reg x_reg_22__retimed_I4062_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4062_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10];
	end
assign N6930 = x_reg_22__retimed_I4062_QOUT;
reg x_reg_22__retimed_I4034_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4034_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638;
	end
assign N6860 = x_reg_22__retimed_I4034_QOUT;
reg x_reg_22__retimed_I4004_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4004_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11];
	end
assign N6784 = x_reg_22__retimed_I4004_QOUT;
reg x_reg_22__retimed_I4001_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I4001_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12];
	end
assign N6777 = x_reg_22__retimed_I4001_QOUT;
reg x_reg_22__retimed_I3904_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3904_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13];
	end
assign N6523 = x_reg_22__retimed_I3904_QOUT;
reg x_reg_22__retimed_I3756_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3756_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0];
	end
assign N6147 = x_reg_22__retimed_I3756_QOUT;
reg x_reg_22__retimed_I3753_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3753_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738;
	end
assign N6138 = x_reg_22__retimed_I3753_QOUT;
reg x_reg_22__retimed_I3741_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3741_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746;
	end
assign N6102 = x_reg_22__retimed_I3741_QOUT;
reg x_reg_22__retimed_I3739_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3739_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439;
	end
assign N6095 = x_reg_22__retimed_I3739_QOUT;
reg x_reg_22__retimed_I3738_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3738_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5];
	end
assign N6093 = x_reg_22__retimed_I3738_QOUT;
reg x_reg_22__retimed_I3736_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3736_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6];
	end
assign N6086 = x_reg_22__retimed_I3736_QOUT;
reg x_reg_22__retimed_I3727_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3727_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2];
	end
assign N6057 = x_reg_22__retimed_I3727_QOUT;
reg x_reg_22__retimed_I3726_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3726_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1];
	end
assign N6055 = x_reg_22__retimed_I3726_QOUT;
reg x_reg_22__retimed_I3718_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3718_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707;
	end
assign N6033 = x_reg_22__retimed_I3718_QOUT;
reg x_reg_22__retimed_I3695_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3695_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681;
	end
assign N5974 = x_reg_22__retimed_I3695_QOUT;
reg x_reg_23__retimed_I3594_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3594_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650;
	end
assign N5705 = x_reg_23__retimed_I3594_QOUT;
reg x_reg_7__retimed_I3592_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3592_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912;
	end
assign N5700 = x_reg_7__retimed_I3592_QOUT;
reg x_reg_31__retimed_I3585_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3585_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6;
	end
assign N5616 = x_reg_31__retimed_I3585_QOUT;
reg x_reg_31__retimed_I3584_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3584_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48;
	end
assign N5614 = x_reg_31__retimed_I3584_QOUT;
reg x_reg_23__retimed_I3576_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3576_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12;
	end
assign N5590 = x_reg_23__retimed_I3576_QOUT;
reg x_reg_23__retimed_I3575_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_23__retimed_I3575_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17;
	end
assign N5588 = x_reg_23__retimed_I3575_QOUT;
reg x_reg_22__retimed_I3572_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_22__retimed_I3572_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63;
	end
assign N5572 = x_reg_22__retimed_I3572_QOUT;
reg x_reg_31__retimed_I3477_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3477_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113;
	end
assign N5336 = x_reg_31__retimed_I3477_QOUT;
reg x_reg_31__retimed_I3476_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_31__retimed_I3476_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122;
	end
assign N5334 = x_reg_31__retimed_I3476_QOUT;
reg x_reg_0__retimed_I3449_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_0__retimed_I3449_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0];
	end
assign N5270 = x_reg_0__retimed_I3449_QOUT;
reg x_reg_1__retimed_I3446_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_1__retimed_I3446_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1];
	end
assign N5263 = x_reg_1__retimed_I3446_QOUT;
reg x_reg_2__retimed_I3443_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_2__retimed_I3443_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2];
	end
assign N5256 = x_reg_2__retimed_I3443_QOUT;
reg x_reg_3__retimed_I3440_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_3__retimed_I3440_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3];
	end
assign N5249 = x_reg_3__retimed_I3440_QOUT;
reg x_reg_4__retimed_I3437_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_4__retimed_I3437_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4];
	end
assign N5242 = x_reg_4__retimed_I3437_QOUT;
reg x_reg_5__retimed_I3434_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_5__retimed_I3434_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5];
	end
assign N5235 = x_reg_5__retimed_I3434_QOUT;
reg x_reg_6__retimed_I3431_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_6__retimed_I3431_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6];
	end
assign N5228 = x_reg_6__retimed_I3431_QOUT;
reg x_reg_7__retimed_I3428_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_7__retimed_I3428_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7];
	end
assign N5221 = x_reg_7__retimed_I3428_QOUT;
reg x_reg_8__retimed_I3425_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_8__retimed_I3425_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8];
	end
assign N5214 = x_reg_8__retimed_I3425_QOUT;
reg x_reg_9__retimed_I3422_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_9__retimed_I3422_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9];
	end
assign N5207 = x_reg_9__retimed_I3422_QOUT;
reg x_reg_10__retimed_I3419_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_10__retimed_I3419_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10];
	end
assign N5200 = x_reg_10__retimed_I3419_QOUT;
reg x_reg_11__retimed_I3416_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_11__retimed_I3416_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11];
	end
assign N5193 = x_reg_11__retimed_I3416_QOUT;
reg x_reg_12__retimed_I3413_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_12__retimed_I3413_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12];
	end
assign N5186 = x_reg_12__retimed_I3413_QOUT;
reg x_reg_13__retimed_I3410_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_13__retimed_I3410_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13];
	end
assign N5179 = x_reg_13__retimed_I3410_QOUT;
reg x_reg_14__retimed_I3407_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_14__retimed_I3407_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14];
	end
assign N5172 = x_reg_14__retimed_I3407_QOUT;
reg x_reg_15__retimed_I3404_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_15__retimed_I3404_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15];
	end
assign N5165 = x_reg_15__retimed_I3404_QOUT;
reg x_reg_16__retimed_I3401_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_16__retimed_I3401_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16];
	end
assign N5158 = x_reg_16__retimed_I3401_QOUT;
reg x_reg_17__retimed_I3398_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_17__retimed_I3398_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17];
	end
assign N5151 = x_reg_17__retimed_I3398_QOUT;
reg x_reg_18__retimed_I3395_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_18__retimed_I3395_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18];
	end
assign N5144 = x_reg_18__retimed_I3395_QOUT;
reg x_reg_19__retimed_I3392_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_19__retimed_I3392_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19];
	end
assign N5137 = x_reg_19__retimed_I3392_QOUT;
reg x_reg_20__retimed_I3389_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_20__retimed_I3389_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20];
	end
assign N5130 = x_reg_20__retimed_I3389_QOUT;
reg x_reg_21__retimed_I3386_QOUT;
always @ (posedge aclk)
	if (bdw_enable==1'b1) begin x_reg_21__retimed_I3386_QOUT <= fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21];
	end
assign N5123 = x_reg_21__retimed_I3386_QOUT;
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I0 (.Y(bdw_enable), .A(astall));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083), .A(a_exp[0]), .B(a_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I2 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085), .A(a_exp[5]), .B(a_exp[4]), .C(a_exp[3]), .D(a_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I3 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194), .A(a_exp[7]), .B(a_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3085));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3083), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8194));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119), .A(a_man[22]), .B(a_man[20]), .C(a_man[21]), .D(a_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I6 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123), .A(a_man[0]), .B(a_man[1]), .C(a_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3119));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I7 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106), .A(a_man[10]), .B(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I8 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125), .A(a_man[6]), .B(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I9 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114), .A(a_man[8]), .B(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I10 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134), .A(a_man[4]), .B(a_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I11 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3106), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3125), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3114), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3134));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I12 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128), .A(a_man[18]), .B(a_man[16]), .C(a_man[17]), .D(a_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I13 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138), .A(a_man[14]), .B(a_man[12]), .C(a_man[13]), .D(a_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I14 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3123), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3117), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3128), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3138));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I15 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I16 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168), .A(b_exp[0]), .B(b_exp[1]));
AND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I17 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170), .A(b_exp[5]), .B(b_exp[4]), .C(b_exp[3]), .D(b_exp[2]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I18 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202), .A(b_exp[7]), .B(b_exp[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3170));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I19 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3168), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8202));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I20 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204), .A(b_man[22]), .B(b_man[20]), .C(b_man[21]), .D(b_man[19]));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I21 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208), .A(b_man[0]), .B(b_man[1]), .C(b_man[2]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3204));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I22 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191), .A(b_man[10]), .B(b_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I23 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210), .A(b_man[6]), .B(b_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I24 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199), .A(b_man[8]), .B(b_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I25 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219), .A(b_man[4]), .B(b_man[3]));
NAND4XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I26 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3210), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3199), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3219));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I27 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213), .A(b_man[18]), .B(b_man[16]), .C(b_man[17]), .D(b_man[15]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I28 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223), .A(b_man[14]), .B(b_man[12]), .C(b_man[13]), .D(b_man[11]));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I29 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3208), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3202), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3213), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3223));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I30 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I31 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__14), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__15));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I32 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__9), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__10));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I33 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]), .A(a_sign), .B(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I34 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I35 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N547));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I36 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .A(b_exp[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I37 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .A(b_exp[6]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I38 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .A(b_exp[5]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I39 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .A(b_exp[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I40 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .A(b_exp[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I41 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .A(b_exp[2]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I42 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .A(b_exp[1]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I43 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .A(b_exp[0]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I44 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I45 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8056));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I46 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3333));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I47 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3327));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I48 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3348));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I49 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3319));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I50 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3343));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I51 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13816));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I52 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13806));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I53 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13813));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I54 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457), .A(a_man[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I55 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .A(b_man[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I56 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544), .A(a_man[21]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I57 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I58 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478), .A(a_man[20]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I59 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I60 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3479));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I61 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3505));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I62 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410), .A(a_man[19]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I63 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I64 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498), .A(a_man[18]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I65 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I66 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I67 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431), .A(a_man[17]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I68 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I69 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515), .A(a_man[16]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I70 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I71 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3537));
NAND3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I72 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3487));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I73 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489), .A(a_man[11]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I74 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I75 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421), .A(a_man[10]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I76 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I77 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3550));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I78 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507), .A(a_man[9]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I79 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I80 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453), .A(a_man[15]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I81 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I82 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535), .A(a_man[14]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I83 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I84 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3492));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I85 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468), .A(a_man[13]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I86 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I87 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405), .A(a_man[12]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I88 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I89 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3446));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I90 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3467));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I91 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444), .A(a_man[8]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I92 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444));
NOR4BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I93 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3503));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I94 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525), .A(a_man[7]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I95 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I96 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461), .A(a_man[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I97 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I98 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3455));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I99 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547), .A(a_man[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I100 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I101 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480), .A(a_man[4]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I102 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I103 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3408));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I104 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3428));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I105 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415), .A(a_man[3]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I106 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I107 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501), .A(a_man[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I108 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I109 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3512));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I110 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441), .A(b_man[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I111 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434), .A(a_man[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I112 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I113 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449), .A(b_man[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3434));
OAI31X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I114 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3441), .A1(a_man[0]), .A2(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3414), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3449));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I115 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546), .A(b_man[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3501));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I116 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494), .A(b_man[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3415));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I117 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3460), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3546), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3494));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I118 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3495), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3527), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3462));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I119 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443), .A(b_man[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3480));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I120 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540), .A(b_man[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3547));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I121 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3506), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3443), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3540));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I122 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488), .A(b_man[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3461));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I123 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437), .A(b_man[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3525));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I124 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3404), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3488), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3437));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I125 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3513), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3548), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3482));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I126 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3504), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3536), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3470));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I127 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534), .A(b_man[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3444));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I128 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483), .A(b_man[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3507));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I129 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3451), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3534), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3483));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I130 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430), .A(b_man[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3421));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I131 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528), .A(b_man[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3489));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I132 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3496), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3430), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3528));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I133 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3532), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3416), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3502));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I134 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477), .A(b_man[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3405));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I135 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424), .A(b_man[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3468));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I136 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3542), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3477), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3424));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I137 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524), .A(b_man[14]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3535));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I138 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471), .A(b_man[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3453));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I139 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3439), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3524), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3471));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I140 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3403), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3436), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3520));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I141 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3522), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3406), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3490));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I142 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3551), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3432), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3517));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I143 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419), .A(b_man[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3515));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I144 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518), .A(b_man[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3431));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I145 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3485), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3419), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3518));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I146 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465), .A(b_man[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3498));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I147 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413), .A(b_man[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3410));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I148 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3530), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3465), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3413));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I149 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3420), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3454), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3539));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I150 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511), .A(b_man[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3478));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I151 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459), .A(b_man[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3544));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I152 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3426), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3511), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3459));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I153 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3475), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3473), .B0(b_man[22]), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3457));
OA21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I154 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3541), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3423), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3508));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I155 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3447), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3499), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3412));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I156 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .A(a_exp[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I157 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N557), .B(a_exp[1]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3321));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I158 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N558), .B(a_exp[2]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3364));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I159 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N559), .B(a_exp[3]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3338));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I160 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N560), .B(a_exp[4]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3358));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I161 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N561), .B(a_exp[5]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3331));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I162 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N562), .B(a_exp[6]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3352));
ADDFX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I163 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N563), .B(a_exp[7]), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3324));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I164 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__34), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I165 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N575));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I166 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I167 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I168 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I169 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .A(a_man[7]), .B(b_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I170 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I171 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269), .A(a_exp[0]), .B(a_exp[7]), .C(a_exp[1]), .D(a_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I172 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273), .A(a_exp[5]), .B(a_exp[3]), .C(a_exp[4]), .D(a_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I173 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3269), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3273));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I174 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291), .A(b_exp[0]), .B(b_exp[7]), .C(b_exp[1]), .D(b_exp[6]));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I175 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295), .A(b_exp[5]), .B(b_exp[3]), .C(b_exp[4]), .D(b_exp[2]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I176 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3291), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3295));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I177 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I178 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I179 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I180 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3701), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N572), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I181 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[1]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I182 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3691), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N566), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I183 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[2]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I184 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3698), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N567), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I185 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I186 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3678), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N569), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I187 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I188 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3671), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N568), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
OAI211X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I189 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]), .C0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I190 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I191 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3694), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N571), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I192 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I193 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3686), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N570), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
NOR3BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I194 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3730), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[6]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[5]));
NAND2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I195 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3729));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I196 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I197 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I198 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N556), .B(a_exp[0]));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I199 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3682), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3688), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N565), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[8]));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I200 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[0]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I201 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I202 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I203 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[1]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I204 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I205 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I206 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__35[4]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I207 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I208 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .A(b_man[12]), .B(a_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I209 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828), .A(b_man[11]), .B(a_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I210 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13828));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I211 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I212 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I213 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .A(b_man[8]), .B(a_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I214 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .A(b_man[7]), .B(a_man[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I215 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I216 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I217 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835), .A(b_man[14]), .B(a_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I218 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13835));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I219 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842), .A(b_man[13]), .B(a_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I220 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13842));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I221 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I222 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .A(b_man[10]), .B(a_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I223 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .A(b_man[9]), .B(a_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I224 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I225 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I226 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I227 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I228 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .A(b_man[20]), .B(a_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I229 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .A(b_man[19]), .B(a_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I230 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I231 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .A(b_man[16]), .B(a_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I232 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .A(b_man[15]), .B(a_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I233 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I234 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I235 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .A(b_man[22]), .B(a_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I236 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .A(b_man[21]), .B(a_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I237 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I238 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .A(b_man[18]), .B(a_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I239 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .A(b_man[17]), .B(a_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I240 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I241 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I242 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I243 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I244 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I245 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I246 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[33]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I247 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8229));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I248 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I249 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .A(a_man[6]), .B(b_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I250 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I251 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I252 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I253 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[37]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[36]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I254 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .A(b_man[6]), .B(a_man[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I255 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[33]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I256 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I257 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[38]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I258 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[34]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I259 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I260 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I261 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I262 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[44]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I263 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[41]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[40]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I264 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I265 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[46]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I266 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[42]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I267 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I268 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I269 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I270 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I271 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[32]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I272 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8222));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I273 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I274 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I275 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3896), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I276 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3960), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I277 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .A(b_man[5]), .B(a_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I278 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[32]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I279 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3979), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I280 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3932));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I281 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I282 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3950), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3926), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I283 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3874));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I284 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I285 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I286 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[31]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I287 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I288 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I289 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629), .A(a_man[5]), .B(b_man[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
AOI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I290 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13607), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13615), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I291 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13597), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13617));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I292 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13629), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13593));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I293 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .A(a_man[4]), .B(b_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I294 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3849));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I295 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3868), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I296 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058), .A(b_man[4]), .B(a_man[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I297 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13058));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I298 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[31]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I299 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3935), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I300 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3881));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I301 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I302 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3877), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3907), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I303 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4044));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I304 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I305 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I306 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[30]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I307 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[30]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I308 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I309 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I310 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4017));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I311 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3986), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I312 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849), .A(b_man[3]), .B(a_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I313 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13849));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I314 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[30]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I315 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3884), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I316 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4053));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I317 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I318 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4047), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3858), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I319 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3996), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I320 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I321 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I322 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[29]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I323 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I324 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .A(a_man[3]), .B(b_man[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13149));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I325 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I326 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I327 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I328 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3942), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3971));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I329 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3893));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I330 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .A(b_man[2]), .B(a_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I331 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[29]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I332 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4056), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I333 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4003));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I334 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I335 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3999), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4027));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I336 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3947));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I337 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I338 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I339 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I340 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I341 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385));
OR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I342 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13376), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13369));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I343 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366), .A(a_man[1]), .B(b_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I344 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4024), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3904));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I345 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I346 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3846), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3968));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I347 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .A(b_man[1]), .B(a_man[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I348 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[28]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I349 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4006), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I350 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3956));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I351 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I352 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I353 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[27]));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I354 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8208));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I355 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I356 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13366));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I357 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I358 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I359 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .A(a_man[0]), .B(b_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I360 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I361 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3923), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4014));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I362 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .A(b_man[0]), .B(a_man[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3769));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I363 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[27]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I364 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3959), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I365 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3911));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I366 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I367 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3975), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3855));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I368 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I369 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I370 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[26]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I371 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13864), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[26]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I372 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
XOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I373 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N655), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I374 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[26]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4021));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I375 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3851), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3915));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I376 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3864));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I377 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3998));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I378 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4042), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I379 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[25]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I380 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[25]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I381 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3867));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I382 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4031));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I383 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3949), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I384 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3994), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I385 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I386 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3883));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I387 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3930));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I388 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3913));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I389 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3985));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I390 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3889), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I391 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3857), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I392 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I393 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3892));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I394 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I395 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I396 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3984));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I397 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4035), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I398 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3901), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4033));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I399 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3983));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I400 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I401 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3958));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I402 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3980), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I403 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I404 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4040), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4041), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4011));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I405 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I406 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3866));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I407 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4008), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I408 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3891));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I409 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4055));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I410 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I411 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[9]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I412 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4363), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4372));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I413 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[14]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4335));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I414 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3934), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3852), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I415 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3928), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I416 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4005));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I417 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4051));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I418 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4012), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3906));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I419 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3869), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I420 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3921), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4026));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I421 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3899));
NOR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I422 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[16]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[15]), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[13]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I423 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4339), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4342));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I424 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4001), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3945), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I425 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3954), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3902));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I426 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3843));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I427 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3962));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I428 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3965), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I429 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3886), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3990));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I430 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[8]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I431 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3919), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3992));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I432 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I433 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4032));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I434 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3916), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I435 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3939));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I436 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3937));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I437 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[10]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I438 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4337), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4346));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I439 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4349));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I440 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3964), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3977), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3993), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I441 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4022), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I442 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3853), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3909));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I443 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4019), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3862));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I444 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3840), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3879));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I445 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[17]));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I446 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3860));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I447 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I448 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I449 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3952), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4049));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I450 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13856), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13858));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I451 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4333), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4343));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I452 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4029), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3973));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I453 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4354), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[19]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I454 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4366), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4351));
NOR3X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I455 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[21]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4356));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I456 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4362), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4332));
AOI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I457 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4353), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4371), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__31));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I458 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I459 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I460 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I461 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13372), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13365), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13389));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I462 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384), .A(a_man[2]), .B(b_man[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13150));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I463 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13385), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13371));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I464 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13384), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13367));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I465 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13354), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I466 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13392), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13387));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I467 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N658), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[4]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I468 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I469 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13608));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I470 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13610));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I471 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13596), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I472 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13635));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I473 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13621), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13601));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I474 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13606));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I475 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N661), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[7]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I476 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4719));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I477 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N662), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[8]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I478 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4647));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I479 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I480 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .A(a_man[8]), .B(b_man[8]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I481 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4046));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I482 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3872), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I483 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[34]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I484 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[34]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I485 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I486 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I487 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4718), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4713));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I488 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I489 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4643), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4648));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I490 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13627));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I491 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13613), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13634), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13611));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I492 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4635), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4586));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I493 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I494 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864));
INVXL buf1_A_I5091 (.Y(N9459), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13599));
INVXL buf1_A_I5092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667), .A(N9459));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I496 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13604));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I497 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4691), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4668));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I498 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4604));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I499 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I500 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13350));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I501 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13378));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I502 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13362));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I503 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4684));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I504 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13388));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I505 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13872));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I506 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13375));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I507 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13877));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I508 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13352));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I509 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13380), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13359));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I510 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4657), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4621));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I511 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I512 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I513 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4845), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I514 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I515 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .A(a_man[15]), .B(b_man[15]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I516 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4037), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I517 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3885), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I518 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[41]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I519 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8250));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I520 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4636), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I521 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .A(a_man[14]), .B(b_man[14]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I522 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3895), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I523 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4007), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I524 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[40]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I525 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[40]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I526 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I527 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .A(a_man[13]), .B(b_man[13]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I528 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3848), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I529 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3914), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I530 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[39]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I531 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[39]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I532 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I533 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .A(a_man[12]), .B(b_man[12]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I534 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4016), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I535 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4034), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I536 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[38]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I537 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[38]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I538 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I539 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .A(a_man[11]), .B(b_man[11]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I540 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3970));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I541 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3940), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I542 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[37]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I543 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8243));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I544 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I545 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .A(a_man[10]), .B(b_man[10]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I546 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3925), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I547 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3844), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I548 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[36]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I549 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8236));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I550 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I551 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .A(a_man[9]), .B(b_man[9]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13148));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I552 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3876), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3920));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I553 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3842), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3966), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I554 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[35]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I555 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[35]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I556 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I557 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N663), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[9]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I558 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4628), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4709), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4579));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I559 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N664), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[10]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I560 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4653));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I561 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N665), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I562 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4589));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I563 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N666), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I564 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4663));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I565 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N667), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I566 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4595));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I567 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N668), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I568 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4673));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I569 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N669), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[15]));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I570 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4659), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4722), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4664), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4603));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I571 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4679), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N670), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[16]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I573 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .A(a_man[16]), .B(b_man[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I574 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3978));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I575 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[42]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I576 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4700), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
DLY1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4961 (.Y(N9213), .A(N8003));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4962 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723), .A0N(N9213), .A1N(N8005), .B0(N8086));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I577 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .A(N7997), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I580 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .A(N8011), .B(N8013));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I581 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4585), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4654));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I584 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4717), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4593));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I585 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4616), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4676));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I586 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I587 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4583), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4610));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I588 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4612), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4692));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I589 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I592 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13145));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I593 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .A(a_man[19]), .B(b_man[19]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I594 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4048));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I595 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[45]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I596 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I597 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .A(a_man[18]), .B(b_man[18]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I598 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3951));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I599 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[44]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I600 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[44]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I601 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4682), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I602 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .A(a_man[17]), .B(b_man[17]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13147));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I603 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3859));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I604 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[43]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I605 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[43]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I606 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4620), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I607 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4609), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N671), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[17]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I609 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4687), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N672), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[18]));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4960 (.Y(N9205), .A(N8003), .B(N8005));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4963 (.Y(N9206), .A(N7997));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4964 (.Y(N9217), .A0(N8086), .A1(N9205), .B0(N9206));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699), .A0N(N7997), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4723), .B0(N8078));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4966 (.Y(N9208), .A(N8078));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I611 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4618), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N673), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[19]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I613 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4695), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N674), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[20]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I615 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .A(a_man[20]), .B(b_man[20]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I616 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3927));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I617 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[46]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I618 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4665), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5049 (.Y(N9361), .A0(N9208), .A1(N9217), .B0(N7990));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5050 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .A(N8070), .B(N9361));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5053 (.Y(N9238), .A0N(N7983), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B0(N8062));
INVXL buf1_A_I5093 (.Y(N9464), .A(N9238));
INVXL buf1_A_I5094 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .A(N9464));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4974 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .A0N(N7976), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .B0(N8054));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I619 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .B(N7969));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I622 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B(N7983));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I623 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4699), .B(N7990));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I626 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .A(a_man[21]), .B(b_man[21]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I627 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4018));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I628 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[47]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I629 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4582), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I630 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N675), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[21]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I632 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4704), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N676), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[22]));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5051 (.Y(N9349), .A(N8062));
AOI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5052 (.Y(N9347), .A0(N7983), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4597), .B0(N9349));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5054 (.Y(N9355), .A(N8054));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5055 (.Y(N9354), .A(N7976));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5056 (.Y(N9348), .A(N9354), .B(N9347));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5057 (.Y(N9236), .A(N9355), .B(N9348));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4975 (.Y(N9239), .A(N7969));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4977 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666), .A0N(N7969), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4578), .B0(N8046));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5085 (.Y(N9448), .A(N8046));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5086 (.Y(N9445), .A(N9239), .B(N9236));
OAI21X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5087 (.Y(N9438), .A0(N9448), .A1(N9445), .B0(N7962));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5088 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672), .A(N8038), .B(N9438));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5089 (.Y(N9441), .A(N7955), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5090 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594), .A(N8030), .B(N9441));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I634 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .A(a_man[22]), .B(b_man[22]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13146));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I635 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3897));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I636 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[48]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I637 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4644), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I638 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4672), .B(N7955));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I639 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .A(N7962), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4666));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I641 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4277), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3890), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3988));
CLKXOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I642 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4677), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4400), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[49]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I643 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8257), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N677), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[23]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I645 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624), .A(N7941), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594));
XOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I646 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]), .A(N7946), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4624));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4983 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .A(N7871), .B(N7873));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5061 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .B(N8148));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5059 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A(N8003), .B(N8005));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5060 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5073 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4984 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5062 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4701), .B(N7976));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5063 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5064 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5065 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5066 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5067 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A(N7941), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4594));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5068 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]));
NAND2X8 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5069 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5070 (.Y(N9387), .AN(N8148), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5071 (.Y(N9397), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5072 (.Y(N9407), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .A1(N9387), .B0(N9397));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5074 (.Y(N9373), .A0(N7820), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826), .B0(N9407));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5075 (.Y(N9381), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5076 (.Y(N9391), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5077 (.Y(N9401), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .A1(N9381), .B0(N9391));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5078 (.Y(N9410), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5079 (.Y(N9377), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]));
OAI21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5080 (.Y(N9385), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A1(N9410), .B0(N9377));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5081 (.Y(N9395), .A0(N9401), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855), .B0(N9385));
NOR2X8 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5082 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855));
AOI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5083 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .A1(N9373), .B0(N9395));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I651 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I652 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I653 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4855));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I654 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4836), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4873), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4893));
OA21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I655 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .A0(N7608), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4913));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I656 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N3367));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I657 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13916));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I658 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I659 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]), .A(a_exp[1]), .B(b_exp[1]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I660 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[2]), .A(a_exp[2]), .B(b_exp[2]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I661 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729), .A(N6055), .B(N6057));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I662 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4837), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4856));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I663 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4896), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4864), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4904), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4883));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I664 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4840), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4894), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4914));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I665 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4850));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I666 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4829), .A1(N7768), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4859));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I667 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4857), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4878));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I668 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4907));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I669 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4885), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4868), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4887));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I670 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4880), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4909));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I671 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .A1(N7662), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4862));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I672 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I674 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5738), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I675 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4872));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I676 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__44), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[0]));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I677 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4639), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4707));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I678 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I679 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[3]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I680 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[5]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I681 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[4]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4869), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4888));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I682 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[7]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I683 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[9]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I684 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[8]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4898), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4918));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I685 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4891), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4910), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4846));
AOI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I686 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4863), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4831), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4848), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4835));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I687 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[11]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I688 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[13]));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I689 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4874), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[12]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4832), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4852));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I702 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]), .A0(N7752), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4905));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I703 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[0]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4876 (.Y(N9073), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4877 (.Y(N9074), .A(N9073));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I704 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .A(a_exp[0]), .B(b_exp[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I705 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I707 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I708 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13151));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I709 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4827), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[0]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I710 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870), .A(N8535), .B(N8533));
NAND2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I711 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I712 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4986 (.Y(N9261), .A(N8533));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4987 (.Y(N9267), .A(N8535), .B(N9261));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4988 (.Y(N9269), .AN(N8535), .B(N8533));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4989 (.Y(N9273), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4892));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4990 (.Y(N9265), .A(N9267), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4900), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4826));
AO21X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4991 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4842), .A1(N9269), .B0(N9273));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4992 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174), .A(N9265), .B(N9273));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I717 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I718 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .B(N7303));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I719 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4846 (.Y(N9015), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4847 (.Y(N9016), .A(N9015));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I720 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288), .A(N6784), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[19]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I721 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5288), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
CLKAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I722 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285), .A(N7364), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I723 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251), .A(N6930), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[18]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I724 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5251), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
INVX12 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I725 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I726 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I727 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I728 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(N7165));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I729 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[23]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I730 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5267), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I731 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(N7343));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I732 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231), .A(N8148), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[22]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I733 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5231), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I734 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I736 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214), .A(N7371), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I737 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217), .A(N6937), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[17]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I738 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5217), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
CLKAND2X3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I739 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143), .A(N7379), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I740 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180), .A(N7172), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I741 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5180), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I742 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I743 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179), .B(N7350));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I744 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196), .A(N6523), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[21]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I745 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5196), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I746 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8180), .B(N7357));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I747 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159), .A(N6777), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[20]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I748 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5159), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I749 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I753 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5275), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5239), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I754 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223), .A(N7379), .B(N7172), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8179));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I755 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[16]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .S0(N9016));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I756 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5178), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5138), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I757 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5254), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5220), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I759 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5205), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5168), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I760 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5183), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5149), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I763 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146), .A(N7165), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[15]), .S0(N9016));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I764 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5146), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I765 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272), .A(N7343), .B(N8148), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I766 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5272));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I767 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5253), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5029 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I770 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5131), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5226), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5030 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I773 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236), .A(N7350), .B(N6523), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8177));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I774 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5236));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I775 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8174));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I776 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202), .A(N7357), .B(N6777), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I777 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5202));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I778 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5031 (.Y(N9298), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5274));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5032 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468));
BUFX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5033 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13468));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5034 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .A0(N9298), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I781 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5155), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5245), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5035 (.Y(N9314), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5036 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(N9314), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I784 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165), .A(N7303), .B(N6784), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I785 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5165), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I786 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5175), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I787 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I788 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5238));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5037 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(N9314), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I790 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128), .A(N7364), .B(N6930), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I791 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5128));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I792 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5266), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I793 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5204));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5038 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .A0(N9298), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5039 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I796 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258), .A(N7371), .B(N6937), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8178));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I797 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5258));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I798 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5223));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I799 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I800 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5129));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I801 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13489));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I802 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13469));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I803 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5162));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I804 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5195), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5287), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I805 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13535), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5166));
OAI2BB1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I806 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13499));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I807 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13513));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I808 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5199));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I809 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I821 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5172), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I822 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5263), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I823 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I813 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I814 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13889));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I824 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13486));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I810 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5152), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I811 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5242), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I812 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I815 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13518), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I825 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I826 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5235), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5164), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I827 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13504));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I817 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5216), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5145), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I818 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13475), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13533));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I828 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I829 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5192), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I830 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5285), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I831 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I832 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5243), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I833 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13540), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I834 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5257), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I835 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5279));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I836 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13483), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I837 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I838 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13503));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I839 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13479));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I816 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13485), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13500));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I819 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13528), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13515));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I820 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
NOR3X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5040 (.Y(N9318), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13478), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13493), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13519));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I841 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5214));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I842 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5143));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I843 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13152), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I844 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5174), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I845 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5206), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I846 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5247), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5278), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5208), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I847 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5210), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I848 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5240), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
NOR2X8 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I849 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5134), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5283));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I850 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5137));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I851 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5169), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I852 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I853 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5132), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I854 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I855 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5265));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I856 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193));
MXI2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I857 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13294), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13298), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I858 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5229));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I859 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5261));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I860 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I873 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13284));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I874 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I875 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .A(N7421), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[0]));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I876 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N631), .B(N7323), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I877 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280), .A(N6860), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I878 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5193));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I879 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211));
MXI2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I880 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[1]), .B(N6953), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I883 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I884 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__54));
CLKAND2X3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I885 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633), .A(N7046), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N632));
NOR4X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I886 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269), .A(N6943), .B(N6945), .C(N6947), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N633));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I887 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269));
MXI2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I888 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5139), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13272), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
OAI21X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I889 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13312), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13275));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I890 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13268), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13305), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13314));
NAND4X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I891 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
INVX3 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5041 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8072));
INVXL buf1_A_I5095 (.Y(N9469), .A(N9318));
INVXL buf1_A_I5096 (.Y(N9303), .A(N9469));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5043 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596), .A(N9303), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5044 (.Y(N9326), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5045 (.Y(N9294), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
NAND2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5046 (.Y(N9312), .A(N9318), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
NOR3X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I5047 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543), .A(N9326), .B(N9294), .C(N9312));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I769 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5141), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4926 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5148), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5290), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I772 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5177), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I861 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .AN(rm[0]), .B(rm[2]), .C(rm[1]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I862 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .A(b_sign), .B(a_sign), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__32));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I863 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I864 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .AN(rm[1]), .B(rm[2]), .C(rm[0]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I865 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I866 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N638), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I867 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I868 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I869 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N626), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30));
AO21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I870 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__30), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N628), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N627));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I871 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N630), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[25]));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I872 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5486), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__43), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__42));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I881 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .AN(rm[2]), .B(rm[1]), .C(rm[0]));
NOR3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I882 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .A(rm[1]), .B(rm[2]), .C(rm[0]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4921 (.Y(N9086), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5181), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5161), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4924 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .A0(N9086), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5213));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4925 (.Y(N9082), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5228), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5218), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5198), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4927 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .A0(N9082), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5171), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5248));
NAND3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4928 (.Y(N9100), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543));
DLY1X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4929 (.Y(N9088), .A(N9100));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4930 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564), .A(N9088));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4931 (.Y(N9101), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]));
NOR2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]), .A(N9101), .B(N9100));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I903 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .A(a_exp[4]), .B(b_exp[4]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I904 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .A(a_exp[3]), .B(b_exp[3]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I905 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754), .A(N8544), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5743));
ADDHX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I906 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .A(N8522), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5716));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I909 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]), .A(a_exp[5]), .B(b_exp[5]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N574));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I910 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5746), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I912 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .A(b_exp[6]), .B(a_exp[6]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I913 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13439), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I917 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .A(b_exp[7]), .B(a_exp[7]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13433));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I918 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742), .A(N8527));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I919 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446), .A(N8527));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4934 (.CO(N9158), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .A(N9074), .B(N6147), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4935 (.CO(N9125), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135), .B(N6138), .CI(N9158));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4936 (.CO(N9151), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5191), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5729), .CI(N9125));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4937 (.CO(N9117), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5754), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5270), .CI(N9151));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4938 (.CO(N9144), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5142), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5724), .CI(N9117));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4939 (.CO(N9168), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5736), .B(N6102), .CI(N9144));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4940 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .A(N6095), .B(N6093), .CI(N9168));
ADDFHXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I920 (.CO(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734), .S(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13446), .B(N6086), .CI(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13697));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I921 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I922 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I927 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I928 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13681), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__17), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__12), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I930 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[7]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I931 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5708));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I932 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13707), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__29[3]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5707));
AO21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I933 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[24]), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[23]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[25]));
NAND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I934 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754), .A(N6055), .B(N6057), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N642));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4941 (.Y(N9121), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4942 (.Y(N9149), .A(N9121));
NOR3X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4943 (.Y(N9115), .A(N9149), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4944 (.Y(N9132), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4945 (.Y(N9136), .A(N9132));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4946 (.Y(N9163), .A(N9136), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]));
INVX2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4947 (.Y(N9172), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13683));
NAND2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4948 (.Y(N9130), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13742), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13710));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4870), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N4841));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .A(N6033), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13754));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4951 (.Y(N9135), .A(N8527), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13734));
NOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4952 (.Y(N9128), .A(N5974), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]));
NOR2X2 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4953 (.Y(N9147), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .B(N9135));
NAND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4954 (.Y(N9156), .A(N9163), .B(N9115));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4955 (.Y(N9127), .A(N9172), .B(N9130));
NOR3X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4956 (.Y(N9161), .A(N9156), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686), .C(N9127));
NAND2X4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4957 (.Y(N9123), .A(N9128), .B(N9147));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I4958 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875), .A(N9123), .B(N9161));
INVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I940 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
CLKINVX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I941 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NOR2BX4 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I942 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .AN(N5572), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I943 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893), .A(rm[0]), .B(rm[1]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I944 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .A(rm[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5893));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I945 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__48), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__5));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I946 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__7), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N652));
NOR3BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I947 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5912), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N653), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4));
AND2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I948 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62), .B(N5700));
NOR2X6 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I949 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .A(N5572), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I950 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I951 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I952 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5575), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[24]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I953 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[22]));
NAND2BXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I954 (.Y(x[22]), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5982));
NOR2BX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I955 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .AN(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I956 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[21]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[21]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[21]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I957 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5564), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[23]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I958 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[21]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I959 (.Y(x[21]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5123), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5939));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I960 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[20]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[20]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[20]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I961 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I962 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8098), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[22]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I963 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[20]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I964 (.Y(x[20]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5130), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5995));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I965 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[19]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[19]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[19]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I966 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5543), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[21]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I967 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[19]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I968 (.Y(x[19]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5137), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5953));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I969 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[18]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[18]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[18]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I970 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5595), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I971 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I972 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5553), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[20]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I973 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8184), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[18]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I974 (.Y(x[18]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5144), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6008));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I975 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[17]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[17]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[17]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I976 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I977 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5591), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[19]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I978 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[17]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I979 (.Y(x[17]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5151), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5966));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I980 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[16]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[16]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[16]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I981 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I982 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5579), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[18]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I983 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[16]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I984 (.Y(x[16]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5158), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5923));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I985 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[15]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[15]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[15]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I986 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5596), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[17]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I987 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[15]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I988 (.Y(x[15]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5165), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5978));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I989 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[14]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[14]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[14]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I990 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13472));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I991 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13904));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I992 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13512));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I993 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13899));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I994 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13523));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I995 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13894));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I996 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I997 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I998 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5580), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I999 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1000 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1001 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5532), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[16]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1002 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[14]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1003 (.Y(x[14]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5172), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5934));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1004 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[13]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[13]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[13]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1005 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5542), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[15]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1006 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8185), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[13]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1007 (.Y(x[13]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5179), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5990));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1008 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[12]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[12]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[12]));
INVXL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1009 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8183));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1010 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1011 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5556), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[14]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1012 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[12]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1013 (.Y(x[12]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5186), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5947));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1014 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[11]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[11]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[11]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1015 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5568), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[13]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1016 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[11]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1017 (.Y(x[11]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5193), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6003));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1018 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[10]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[10]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[10]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1019 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5539), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1020 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1021 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5583), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[12]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1022 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[10]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1023 (.Y(x[10]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5200), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5961));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1024 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[9]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[9]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[9]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1025 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5567), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[11]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1026 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[9]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1027 (.Y(x[9]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5207), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5918));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1028 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[8]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[8]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[8]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1029 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1030 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8092), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[10]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1031 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8186), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[8]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1032 (.Y(x[8]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5214), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5973));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1033 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[7]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[7]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[7]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1034 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5588), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[9]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1035 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[7]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1036 (.Y(x[7]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5221), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5930));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1037 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[6]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[6]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[6]));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1038 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5546), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1039 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1040 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5561), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[8]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1041 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[6]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1042 (.Y(x[6]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5228), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5986));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1043 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[5]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[5]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[5]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1044 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5594), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[7]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1045 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[5]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1046 (.Y(x[5]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5235), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5943));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1047 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[4]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[4]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[4]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1048 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1049 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5587), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[6]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1050 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[4]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1051 (.Y(x[4]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5242), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5999));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1052 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[3]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[3]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1053 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5557), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[5]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1054 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[3]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1055 (.Y(x[3]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5249), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5956));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1056 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[2]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[2]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[2]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1057 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5211), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5189), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5135));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1058 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13269), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13309));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1059 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13908), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13280));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1060 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]));
NAND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1061 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600));
XNOR2X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1062 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5538), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[4]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1063 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[2]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1064 (.Y(x[2]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5256), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N6011));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1065 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[1]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[1]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[1]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1066 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5600), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[3]));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1067 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[1]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1068 (.Y(x[1]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5263), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5969));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1069 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[0]), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .A1(a_man[0]), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_man[0]));
XOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1070 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__50[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__55));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1071 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__70), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5997), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N8188), .B1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__57[0]));
OAI2BB1XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1072 (.Y(x[0]), .A0N(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5942), .A1N(N5270), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5926));
INVXL buf1_A_I5097 (.Y(N9474), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13686));
INVXL buf1_A_I5098 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .A(N9474));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1074 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .A(N5590), .B(N5588), .C(N5572), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
INVX1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1075 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5875));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1076 (.Y(x[30]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[7]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1077 (.Y(x[29]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[6]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1078 (.Y(x[28]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[5]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1079 (.Y(x[27]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[4]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1080 (.Y(x[26]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[3]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1081 (.Y(x[25]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[2]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1082 (.Y(x[24]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[1]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5869), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1083 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N650), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__4), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__8), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N635), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N634));
AND2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1084 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651), .A(N5705), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__62));
OR4X1 fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1085 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .A(N5588), .B(N5590), .C(N5572), .D(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N651));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1086 (.Y(x[23]), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[0]), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[0]), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5857));
OR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1087 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881), .A(a_sign), .B(b_sign));
AO22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1088 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N13881), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__6), .B0(a_sign), .B1(b_sign));
AND3XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1089 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__11), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__16), .C(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N645));
AOI22XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1090 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064), .A0(a_sign), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5043), .B1(b_sign));
OAI21XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1091 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .A0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__18), .A1(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__13), .B0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5064));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1092 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5113), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__66), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N710), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1093 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .A(N5614), .B(N5616), .S0(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[5]));
NOR2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1094 (.Y(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5122), .A(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__63), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N706));
MX2XL fp_add_cynw_cm_float_add2_ieee_E8_M23_4_I1095 (.Y(x[31]), .A(N5336), .B(fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_N5116), .S0(N5334));
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__27[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[27] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[28] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[31] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[32] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[33] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[36] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[37] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__33[41] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[0] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[7] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[10] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[11] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[12] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[13] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[14] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[15] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[16] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[17] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[18] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[19] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[20] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[21] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[23] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[25] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__36[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[42] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[45] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[46] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[47] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[48] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__37[49] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__39[24] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__45[26] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__49[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[8] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__59[9] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__64[22] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[1] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[2] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[3] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[4] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[5] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[6] = 1'B0;
assign fp_add_cynw_cm_float_add2_ieee_E8_M23_3_inst_inst_cellmath__68[7] = 1'B0;
endmodule

/* CADENCE  v7L3SQHWqhs= : u9/ySgnWtBlWxVPRXgAZ4Og= ** DO NOT EDIT THIS LINE **/



