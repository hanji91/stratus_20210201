`timescale 1ps / 1ps
module fp_cmp_cynw_cm_float_ltle_4_2(
          in1,
          in2,
          in3,
          in4,
          in5,
          in6,
          out1,
          clk
);
   input in1;
   input [7:0] in2;
   input [22:0] in3;
   input [7:0] in4;
   input [22:0] in5;
   input in6;
   output [1:0] out1;
   input clk;
wire asc021, gt_90_21_n_0, gt_90_21_n_1, gt_90_21_n_2, gt_90_21_n_3,
     gt_90_21_n_4, gt_90_21_n_5, gt_90_21_n_6, gt_90_21_n_7, gt_90_21_n_8,
     gt_90_21_n_9, gt_90_21_n_10, gt_90_21_n_11, gt_90_21_n_12, gt_90_21_n_13,
     gt_90_21_n_14, gt_90_21_n_15, gt_90_21_n_16, gt_90_21_n_17, gt_90_21_n_18,
     gt_90_21_n_19, gt_90_21_n_20, gt_90_21_n_21, gt_92_21_n_0, gt_92_21_n_1,
     gt_92_21_n_2, gt_92_21_n_3, gt_92_21_n_4, gt_92_21_n_5, gt_92_21_n_6,
     gt_92_21_n_7, gt_92_21_n_8, gt_92_21_n_9, gt_92_21_n_10, gt_92_21_n_11,
     gt_92_21_n_12, gt_92_21_n_13, gt_92_21_n_14, gt_92_21_n_15, gt_92_21_n_16,
     gt_92_21_n_17, gt_92_21_n_18, gt_92_21_n_19, gt_92_21_n_20, gt_92_21_n_21,
     gt_94_21_n_0, gt_94_21_n_1, gt_94_21_n_2, gt_94_21_n_3, gt_94_21_n_4,
     gt_94_21_n_5, gt_94_21_n_6, gt_94_21_n_7, gt_94_21_n_8, gt_94_21_n_9,
     gt_94_21_n_10, gt_94_21_n_11, gt_94_21_n_12, gt_94_21_n_13, gt_94_21_n_14,
     gt_94_21_n_15, gt_94_21_n_16, gt_94_21_n_17, gt_94_21_n_18, gt_94_21_n_19,
     gt_94_21_n_20, gt_94_21_n_21, gt_94_21_n_22, gt_94_21_n_23, gt_94_21_n_24,
     gt_94_21_n_25, gt_94_21_n_26, gt_94_21_n_27, gt_94_21_n_28, gt_94_21_n_29,
     gt_94_21_n_31, gt_94_21_n_32, gt_94_21_n_33, gt_94_21_n_34, gt_94_21_n_35,
     gt_94_21_n_36, gt_94_21_n_37, gt_94_21_n_38, gt_94_21_n_39, gt_94_21_n_40,
     gt_94_21_n_41, gt_94_21_n_42, gt_94_21_n_43, gt_94_21_n_44, gt_94_21_n_45,
     gt_94_21_n_46, gt_94_21_n_47, gt_94_21_n_48, gt_94_21_n_49, gt_94_21_n_50,
     gt_94_21_n_51, gt_94_21_n_52, gt_94_21_n_53, gt_94_21_n_54, gt_94_21_n_55,
     gt_94_21_n_56, gt_94_21_n_57, gt_94_21_n_58, gt_94_21_n_59, gt_94_21_n_60,
     gt_94_21_n_61, gt_94_21_n_62, gt_94_21_n_63, gt_94_21_n_64, gt_94_21_n_65,
     gt_94_21_n_66, gt_94_21_n_67, gt_94_21_n_68, gt_96_21_n_5, gt_96_21_n_6,
     gt_96_21_n_7, gt_96_21_n_8, gt_96_21_n_9, gt_96_21_n_11, gt_96_21_n_14,
     gt_96_21_n_15, gt_96_21_n_17, gt_96_21_n_19, gt_96_21_n_22, gt_96_21_n_26,
     gt_96_21_n_27, gt_96_21_n_28, gt_96_21_n_29, gt_96_21_n_33, gt_96_21_n_34,
     gt_96_21_n_35, gt_96_21_n_36, gt_96_21_n_37, gt_96_21_n_38, gt_96_21_n_39,
     gt_96_21_n_48, gt_96_21_n_49, gt_96_21_n_50, gt_96_21_n_56, gt_96_21_n_57,
     gt_96_21_n_66, gt_96_21_n_68, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9,
     n_10, n_11, clk, in6, in1, n_15, n_16, n_17, n_19, n_20, n_21, n_22, n_23,
     n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35,
     n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47,
     n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_59, n_60,
     n_61, n_62, n_63, n_64, n_65, n_66, n_67;
assign {out1[0]} = asc021;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         retime_s1_9_reg_reg_N30 <= n_22;
 assign n_3 = retime_s1_9_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         retime_s1_8_reg_reg_N30 <= n_24;
 assign n_4 = retime_s1_8_reg_reg_N30;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= n_47;
 assign n_11 = retime_s1_1_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         retime_s1_10_reg_reg_N30 <= n_49;
 assign n_2 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         retime_s1_11_reg_reg_N30 <= in1;
 assign n_1 = retime_s1_11_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         retime_s1_7_reg_reg_N30 <= {in2[0]};
 assign n_5 = retime_s1_7_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= n_46;
 assign n_10 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= n_25;
 assign n_9 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= n_15;
 assign n_8 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= n_23;
 assign n_7 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= {in2[1]};
 assign n_6 = retime_s1_6_reg_reg_N30;
 assign asc021 = ~(n_19 | (n_5 & (n_6 & n_9)));
 assign n_19 = ~((n_20 | n_21) & (n_4 | n_2));
 assign n_20 = ~((n_3 & n_41) | (n_7 & n_1));
 assign n_21 = ~(n_11 | (n_8 | (n_3 | n_10)));
 assign n_22 = ~(in6 & ({in4[4]} | ({in4[5]} | n_26)));
 assign n_23 = ~(n_27 & (n_39 & (n_50 & n_53)));
 assign n_24 = ~(n_28 & ({in4[2]} & ({in4[3]} & ~n_38)));
 assign n_25 = ~(n_27 | (n_37 | (~{in2[2]} | ~{in2[3]})));
 assign n_26 = (n_28 | (n_40 | ({in4[6]} | {in4[7]})));
 assign n_27 = ~({in3[19]} | ({in3[20]} | ~n_29));
 assign n_28 = ~(n_31 & (n_43 & (n_54 & n_51)));
 assign n_29 = ~(n_30 | (n_45 | ({in3[21]} | {in3[22]})));
 assign n_30 = ~(n_33 & (n_44 & (n_52 & n_48)));
 assign n_31 = ~(n_32 | (n_55 | ({in5[11]} | {in5[12]})));
 assign n_32 = ~(n_34 & n_42);
 assign n_33 = ~(n_36 | ({in3[3]} | ({in3[4]} | {in3[5]})));
 assign n_34 = ~(n_35 | ({in5[3]} | ({in5[4]} | {in5[5]})));
 assign n_35 = ({in5[1]} | ({in5[2]} | ({in5[0]} | {in5[6]})));
 assign n_36 = ({in3[1]} | ({in3[2]} | ({in3[0]} | {in3[6]})));
 assign n_37 = ~({in2[4]} & ({in2[5]} & ({in2[6]} & {in2[7]})));
 assign n_38 = ~({in4[4]} & ({in4[5]} & ({in4[6]} & {in4[7]})));
 assign n_39 = ~({in2[4]} | ({in2[5]} | ({in2[6]} | {in2[7]})));
 assign n_40 = ({in4[0]} | ({in4[1]} | ({in4[2]} | {in4[3]})));
 assign n_41 = ~(n_11 | n_8);
 assign n_42 = ~({in5[7]} | ({in5[8]} | ({in5[9]} | {in5[10]})));
 assign n_43 = ~({in5[19]} | ({in5[20]} | ({in5[21]} | {in5[22]})));
 assign n_44 = ~({in3[7]} | ({in3[8]} | ({in3[9]} | {in3[10]})));
 assign n_45 = ({in3[15]} | ({in3[16]} | ({in3[17]} | {in3[18]})));
 assign n_46 = ~(n_16 | (n_17 | (n_15 | n_56)));
 assign n_47 = ~(n_16 | ~n_17);
 assign n_48 = ~({in3[11]} | {in3[12]});
 assign n_49 = ~({in4[0]} & {in4[1]});
 assign n_50 = ~({in2[2]} | {in2[3]});
 assign n_51 = ~({in5[15]} | {in5[16]});
 assign n_52 = ~({in3[13]} | {in3[14]});
 assign n_53 = ~({in2[0]} | {in2[1]});
 assign n_54 = ~({in5[17]} | {in5[18]});
 assign n_55 = ({in5[13]} | {in5[14]});
 assign n_15 = ~(gt_90_21_n_21 | gt_90_21_n_19);
 assign gt_90_21_n_21 = ~(gt_90_21_n_20 | (gt_90_21_n_11 | (gt_90_21_n_7 | gt_90_21_n_9)));
 assign gt_90_21_n_20 = ~(gt_90_21_n_18 | ((gt_90_21_n_13 & {in4[2]}) | (gt_90_21_n_5 & {in4[3]})));
 assign gt_90_21_n_19 = ~(gt_90_21_n_15 & (({in2[7]} | gt_90_21_n_4) & (gt_90_21_n_16 | gt_90_21_n_11)));
 assign gt_90_21_n_18 = ~(gt_90_21_n_17 | (gt_90_21_n_10 | (gt_90_21_n_3 & {in2[2]})));
 assign gt_90_21_n_17 = ~((gt_90_21_n_12 & {in4[1]}) | (gt_90_21_n_8 & gt_90_21_n_2));
 assign gt_90_21_n_16 = ~((gt_90_21_n_14 & {in4[4]}) | (gt_90_21_n_1 & {in4[5]}));
 assign gt_90_21_n_15 = ~(gt_90_21_n_6 & ({in4[6]} & ~{in2[6]}));
 assign gt_90_21_n_14 = ~(gt_90_21_n_9 | {in2[4]});
 assign gt_90_21_n_13 = ~(gt_90_21_n_10 | {in2[2]});
 assign gt_90_21_n_12 = ~({in2[0]} & ({in2[1]} & ~{in4[0]}));
 assign gt_90_21_n_11 = ~(gt_90_21_n_6 & ({in4[6]} | gt_90_21_n_0));
 assign gt_90_21_n_10 = ~({in4[3]} | gt_90_21_n_5);
 assign gt_90_21_n_9 = ~({in4[5]} | gt_90_21_n_1);
 assign gt_90_21_n_8 = ~({in2[0]} & ~{in4[0]});
 assign gt_90_21_n_7 = ~({in4[4]} | ~{in2[4]});
 assign gt_90_21_n_6 = ~(gt_90_21_n_4 & {in2[7]});
 assign gt_90_21_n_5 = ~{in2[3]};
 assign gt_90_21_n_4 = ~{in4[7]};
 assign gt_90_21_n_3 = ~{in4[2]};
 assign gt_90_21_n_2 = ~{in2[1]};
 assign gt_90_21_n_1 = ~{in2[5]};
 assign gt_90_21_n_0 = ~{in2[6]};
 assign n_16 = ~(gt_92_21_n_21 | gt_92_21_n_19);
 assign gt_92_21_n_21 = ~(gt_92_21_n_20 | (gt_92_21_n_11 | (gt_92_21_n_7 | gt_92_21_n_9)));
 assign gt_92_21_n_20 = ~(gt_92_21_n_18 | ((gt_92_21_n_13 & {in2[2]}) | (gt_92_21_n_5 & {in2[3]})));
 assign gt_92_21_n_19 = ~(gt_92_21_n_15 & (({in4[7]} | gt_92_21_n_4) & (gt_92_21_n_16 | gt_92_21_n_11)));
 assign gt_92_21_n_18 = ~(gt_92_21_n_17 | (gt_92_21_n_10 | (gt_92_21_n_3 & {in4[2]})));
 assign gt_92_21_n_17 = ~((gt_92_21_n_12 & {in2[1]}) | (gt_92_21_n_8 & gt_92_21_n_2));
 assign gt_92_21_n_16 = ~((gt_92_21_n_14 & {in2[4]}) | (gt_92_21_n_1 & {in2[5]}));
 assign gt_92_21_n_15 = ~(gt_92_21_n_6 & ({in2[6]} & ~{in4[6]}));
 assign gt_92_21_n_14 = ~(gt_92_21_n_9 | {in4[4]});
 assign gt_92_21_n_13 = ~(gt_92_21_n_10 | {in4[2]});
 assign gt_92_21_n_12 = ~({in4[0]} & ({in4[1]} & ~{in2[0]}));
 assign gt_92_21_n_11 = ~(gt_92_21_n_6 & ({in2[6]} | gt_92_21_n_0));
 assign gt_92_21_n_10 = ~({in2[3]} | gt_92_21_n_5);
 assign gt_92_21_n_9 = ~({in2[5]} | gt_92_21_n_1);
 assign gt_92_21_n_8 = ~({in4[0]} & ~{in2[0]});
 assign gt_92_21_n_7 = ~({in2[4]} | ~{in4[4]});
 assign gt_92_21_n_6 = ~(gt_92_21_n_4 & {in4[7]});
 assign gt_92_21_n_5 = ~{in4[3]};
 assign gt_92_21_n_4 = ~{in2[7]};
 assign gt_92_21_n_3 = ~{in2[2]};
 assign gt_92_21_n_2 = ~{in4[1]};
 assign gt_92_21_n_1 = ~{in4[5]};
 assign gt_92_21_n_0 = ~{in4[6]};
 assign n_17 = ~((gt_94_21_n_68 | gt_94_21_n_18) & ({in5[22]} | gt_94_21_n_7));
 assign gt_94_21_n_68 = ~(gt_94_21_n_67 & (gt_94_21_n_45 & ({in3[21]} | gt_94_21_n_2)));
 assign gt_94_21_n_67 = ~(gt_94_21_n_25 & ((gt_94_21_n_66 | gt_94_21_n_60) & ({in5[20]} | gt_94_21_n_6)));
 assign gt_94_21_n_66 = ~(gt_94_21_n_65 | (gt_94_21_n_31 | (gt_94_21_n_39 | gt_94_21_n_27)));
 assign gt_94_21_n_65 = ~(gt_94_21_n_64 | (gt_94_21_n_59 | (gt_94_21_n_61 & gt_94_21_n_51)));
 assign gt_94_21_n_64 = ~(gt_94_21_n_50 | (gt_94_21_n_49 | (gt_94_21_n_63 & gt_94_21_n_58)));
 assign gt_94_21_n_63 = ~(gt_94_21_n_62 & (gt_94_21_n_28 & (gt_94_21_n_34 & gt_94_21_n_22)));
 assign gt_94_21_n_62 = ~(gt_94_21_n_57 & (gt_94_21_n_46 & ({in3[3]} | gt_94_21_n_16)));
 assign gt_94_21_n_61 = ~(gt_94_21_n_47 & (({in3[11]} | gt_94_21_n_10) & (gt_94_21_n_54 | gt_94_21_n_37)));
 assign gt_94_21_n_60 = ~(gt_94_21_n_43 & (({in3[19]} | gt_94_21_n_1) & (gt_94_21_n_55 | gt_94_21_n_39)));
 assign gt_94_21_n_59 = ~(gt_94_21_n_44 & (({in3[15]} | gt_94_21_n_13) & (gt_94_21_n_53 | gt_94_21_n_35)));
 assign gt_94_21_n_58 = ~(n_59 | ((gt_94_21_n_52 & gt_94_21_n_34) | (gt_94_21_n_40 & {in5[6]})));
 assign gt_94_21_n_57 = ~(gt_94_21_n_56 & (gt_94_21_n_32 & ({in5[2]} | gt_94_21_n_17)));
 assign gt_94_21_n_56 = ~(gt_94_21_n_48 & (gt_94_21_n_29 | {in3[1]}));
 assign gt_94_21_n_55 = ~((gt_94_21_n_41 & {in5[16]}) | (gt_94_21_n_4 & {in5[17]}));
 assign gt_94_21_n_54 = ~((gt_94_21_n_33 & (gt_94_21_n_8 & {in5[8]})) | (gt_94_21_n_12 & {in5[9]}));
 assign gt_94_21_n_53 = ~((gt_94_21_n_19 & (gt_94_21_n_11 & {in5[12]})) | (gt_94_21_n_0 & {in5[13]}));
 assign gt_94_21_n_52 = ~(gt_94_21_n_42 & ~(gt_94_21_n_3 & {in5[5]}));
 assign gt_94_21_n_51 = ~gt_94_21_n_50;
 assign gt_94_21_n_50 = ~(gt_94_21_n_36 & (gt_94_21_n_19 & ({in5[12]} | gt_94_21_n_11)));
 assign gt_94_21_n_49 = ~(gt_94_21_n_38 & (gt_94_21_n_33 & ({in5[8]} | gt_94_21_n_8)));
 assign gt_94_21_n_48 = ~({in5[1]} & (gt_94_21_n_26 | {in5[0]}));
 assign gt_94_21_n_47 = ~(gt_94_21_n_21 & ({in5[10]} & ~{in3[10]}));
 assign gt_94_21_n_46 = ~(gt_94_21_n_32 & (gt_94_21_n_17 & {in5[2]}));
 assign gt_94_21_n_45 = ~(gt_94_21_n_25 & ({in5[20]} & ~{in3[20]}));
 assign gt_94_21_n_44 = ~(gt_94_21_n_20 & ({in5[14]} & ~{in3[14]}));
 assign gt_94_21_n_43 = ~(gt_94_21_n_24 & ({in5[18]} & ~{in3[18]}));
 assign gt_94_21_n_42 = ~(gt_94_21_n_22 & ({in5[4]} & ~{in3[4]}));
 assign gt_94_21_n_41 = ~(gt_94_21_n_31 | {in3[16]});
 assign gt_94_21_n_40 = ~(gt_94_21_n_23 | {in3[6]});
 assign gt_94_21_n_39 = ~(gt_94_21_n_24 & ({in5[18]} | gt_94_21_n_9));
 assign gt_94_21_n_38 = ~gt_94_21_n_37;
 assign gt_94_21_n_37 = ~(gt_94_21_n_21 & ~(gt_94_21_n_5 & {in3[10]}));
 assign gt_94_21_n_36 = ~gt_94_21_n_35;
 assign gt_94_21_n_35 = ~(gt_94_21_n_20 & ~(gt_94_21_n_14 & {in3[14]}));
 assign gt_94_21_n_34 = ~(gt_94_21_n_23 | (gt_94_21_n_15 & {in3[6]}));
 assign gt_94_21_n_29 = ~({in5[0]} | ~{in3[0]});
 assign gt_94_21_n_28 = ~({in3[4]} & ~{in5[4]});
 assign gt_94_21_n_27 = ~({in5[16]} | ~{in3[16]});
 assign gt_94_21_n_26 = ~({in3[0]} & {in3[1]});
 assign gt_94_21_n_33 = ~({in3[9]} & ~{in5[9]});
 assign gt_94_21_n_32 = ~(gt_94_21_n_16 & {in3[3]});
 assign gt_94_21_n_31 = ~({in5[17]} | gt_94_21_n_4);
 assign gt_94_21_n_18 = ~({in3[22]} | ~{in5[22]});
 assign gt_94_21_n_25 = ~(gt_94_21_n_2 & {in3[21]});
 assign gt_94_21_n_24 = ~(gt_94_21_n_1 & {in3[19]});
 assign gt_94_21_n_23 = ~({in5[7]} | ~{in3[7]});
 assign gt_94_21_n_22 = ~({in3[5]} & ~{in5[5]});
 assign gt_94_21_n_21 = ~(gt_94_21_n_10 & {in3[11]});
 assign gt_94_21_n_20 = ~(gt_94_21_n_13 & {in3[15]});
 assign gt_94_21_n_19 = ~({in3[13]} & ~{in5[13]});
 assign gt_94_21_n_17 = ~{in3[2]};
 assign gt_94_21_n_16 = ~{in5[3]};
 assign gt_94_21_n_15 = ~{in5[6]};
 assign gt_94_21_n_14 = ~{in5[14]};
 assign gt_94_21_n_13 = ~{in5[15]};
 assign gt_94_21_n_12 = ~{in3[9]};
 assign gt_94_21_n_11 = ~{in3[12]};
 assign gt_94_21_n_10 = ~{in5[11]};
 assign gt_94_21_n_9 = ~{in3[18]};
 assign gt_94_21_n_8 = ~{in3[8]};
 assign gt_94_21_n_7 = ~{in3[22]};
 assign gt_94_21_n_6 = ~{in3[20]};
 assign gt_94_21_n_5 = ~{in5[10]};
 assign gt_94_21_n_4 = ~{in3[17]};
 assign gt_94_21_n_3 = ~{in3[5]};
 assign gt_94_21_n_2 = ~{in5[21]};
 assign gt_94_21_n_1 = ~{in5[19]};
 assign gt_94_21_n_0 = ~{in3[13]};
 assign gt_96_21_n_66 = ~(n_60 | (n_64 | (gt_96_21_n_39 | gt_96_21_n_27)));
 assign gt_96_21_n_57 = ~(gt_96_21_n_56 & (n_61 & ({in3[2]} | gt_96_21_n_17)));
 assign gt_96_21_n_56 = ~(gt_96_21_n_48 & (gt_96_21_n_29 | {in5[1]}));
 assign gt_96_21_n_50 = ~(gt_96_21_n_36 & (gt_96_21_n_19 & ({in3[12]} | gt_96_21_n_11)));
 assign gt_96_21_n_49 = ~(gt_96_21_n_38 & (gt_96_21_n_33 & ({in3[8]} | gt_96_21_n_8)));
 assign gt_96_21_n_48 = ~({in3[1]} & (gt_96_21_n_26 | {in3[0]}));
 assign gt_96_21_n_39 = ~(n_66 & ({in3[18]} | gt_96_21_n_9));
 assign gt_96_21_n_38 = ~gt_96_21_n_37;
 assign gt_96_21_n_37 = ~(n_63 & ~(gt_96_21_n_5 & {in5[10]}));
 assign gt_96_21_n_36 = ~gt_96_21_n_35;
 assign gt_96_21_n_35 = ~(n_62 & ~(gt_96_21_n_14 & {in5[14]}));
 assign gt_96_21_n_34 = ~(n_59 | (gt_96_21_n_15 & {in5[6]}));
 assign gt_96_21_n_29 = ~({in3[0]} | ~{in5[0]});
 assign gt_96_21_n_28 = ~({in5[4]} & ~{in3[4]});
 assign gt_96_21_n_27 = ~({in3[16]} | ~{in5[16]});
 assign gt_96_21_n_33 = ~({in5[9]} & ~{in3[9]});
 assign gt_96_21_n_22 = ~({in5[5]} & ~{in3[5]});
 assign gt_96_21_n_19 = ~({in5[13]} & ~{in3[13]});
 assign gt_96_21_n_17 = ~{in5[2]};
 assign gt_96_21_n_15 = ~{in3[6]};
 assign gt_96_21_n_14 = ~{in3[14]};
 assign gt_96_21_n_11 = ~{in5[12]};
 assign gt_96_21_n_9 = ~{in5[18]};
 assign gt_96_21_n_8 = ~{in5[8]};
 assign gt_96_21_n_7 = ~{in5[22]};
 assign gt_96_21_n_6 = ~{in5[20]};
 assign gt_96_21_n_5 = ~{in3[10]};
 assign gt_96_21_n_26 = ~{in5[0]};
 assign gt_96_21_n_68 = ~n_57;
 assign n_56 = ~(gt_96_21_n_68 & ({in3[22]} | gt_96_21_n_7));
 assign n_57 = ~(n_65 & (gt_96_21_n_66 & ({in3[20]} | gt_96_21_n_6)));
 assign n_59 = ~({in3[7]} | ~{in5[7]});
 assign n_60 = (gt_96_21_n_50 | (gt_96_21_n_49 | n_67));
 assign n_61 = ~({in5[3]} & ~{in3[3]});
 assign n_62 = ~({in5[15]} & ~{in3[15]});
 assign n_63 = ~({in5[11]} & ~{in3[11]});
 assign n_64 = ~({in3[17]} | ~{in5[17]});
 assign n_65 = ~({in5[21]} & ~{in3[21]});
 assign n_66 = ~({in5[19]} & ~{in3[19]});
 assign n_67 = ~(gt_96_21_n_28 & (gt_96_21_n_34 & (gt_96_21_n_22 & ~gt_96_21_n_57)));
assign out1[1] = 1'B0;
endmodule

